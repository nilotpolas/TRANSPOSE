module sbox(
    clk,
    t,
    dec_0,
    dec_1,
    dec_255,
    dec_169,
    dec_129,
    dec_9,
    dec_72,
    dec_242,
    dec_243,
    dec_152,
    dec_240,
    dec_4,
    dec_15,
    dec_12,
    dec_2,
    dec_3,
    dec_36,
    dec_220,
    dec_11,
    dec_158,
    dec_45,
    dec_88,
    dec_99,
    r,
    y
);
//inputS
    input clk;
    input [7:0]  t;
    input [7:0]  dec_0;
    input [7:0]  dec_1;
    input [7:0]  dec_255;
    input [7:0]  dec_169;
    input [7:0]  dec_129;
    input [7:0]  dec_9;
    input [7:0]  dec_72;
    input [7:0]  dec_242;
    input [7:0]  dec_243;
    input [7:0]  dec_152;
    input [7:0]  dec_240;
    input [7:0]  dec_4;
    input [7:0]  dec_15;
    input [7:0]  dec_12;
    input [7:0]  dec_2;
    input [7:0]  dec_3;
    input [7:0]  dec_36;
    input [7:0]  dec_220;
    input [7:0]  dec_11;
    input [7:0]  dec_158;
    input [7:0]  dec_45;
    input [7:0]  dec_88;
    input [7:0]  dec_99;
	input [20:0] r;
//OUTPUTS
    output reg [7:0]  y;
//Intermediate values
    wire [7:0] dec_99_inp;
    wire [7:0] dec_88_inp;
    wire [7:0] dec_45_inp;
    wire [7:0] dec_158_inp;
    wire [7:0] dec_11_inp;
    wire [7:0] dec_220_inp;
    wire [7:0] dec_36_inp;
    wire [7:0] dec_3_inp;
    wire [7:0] dec_2_inp;
    wire [7:0] dec_12_inp;
    wire [7:0] dec_15_inp;
    wire [7:0] dec_4_inp;
    wire [7:0] dec_240_inp;
    wire [7:0] dec_152_inp;
    wire [7:0] dec_243_inp;
    wire [7:0] dec_242_inp;
    wire [7:0] dec_72_inp;
    wire [7:0] dec_9_inp;
    wire [7:0] dec_129_inp;
    wire [7:0] dec_169_inp;
    wire [7:0] dec_255_inp;
    wire [7:0] dec_1_inp;
    wire [7:0] dec_0_inp;
    wire [7:0] t_inp;
    wire [7:0] y_G256_newbasis0;
    wire [7:0] tempy1_G256_newbasis0;
    wire [7:0] cond1_G256_newbasis0;
    wire [7:0] negCond1_G256_newbasis0;
    wire [7:0] yxorb1_G256_newbasis0;
    wire [7:0] ny1_G256_newbasis0;
    wire [7:0] tempyIntoNegCond1_G256_newbasis0;
    wire [7:0] y1_G256_newbasis0;
    wire [7:0] x1_G256_newbasis0;
    wire [7:0] tempy2_G256_newbasis0;
    wire [7:0] cond2_G256_newbasis0;
    wire [7:0] negCond2_G256_newbasis0;
    wire [7:0] yxorb2_G256_newbasis0;
    wire [7:0] ny2_G256_newbasis0;
    wire [7:0] tempyIntoNegCond2_G256_newbasis0;
    wire [7:0] y2_G256_newbasis0;
    wire [7:0] x2_G256_newbasis0;
    wire [7:0] tempy3_G256_newbasis0;
    wire [7:0] cond3_G256_newbasis0;
    wire [7:0] negCond3_G256_newbasis0;
    wire [7:0] yxorb3_G256_newbasis0;
    wire [7:0] ny3_G256_newbasis0;
    wire [7:0] tempyIntoNegCond3_G256_newbasis0;
    wire [7:0] y3_G256_newbasis0;
    wire [7:0] x3_G256_newbasis0;
    wire [7:0] tempy4_G256_newbasis0;
    wire [7:0] cond4_G256_newbasis0;
    wire [7:0] negCond4_G256_newbasis0;
    wire [7:0] yxorb4_G256_newbasis0;
    wire [7:0] ny4_G256_newbasis0;
    wire [7:0] tempyIntoNegCond4_G256_newbasis0;
    wire [7:0] y4_G256_newbasis0;
    wire [7:0] x4_G256_newbasis0;
    wire [7:0] tempy5_G256_newbasis0;
    wire [7:0] cond5_G256_newbasis0;
    wire [7:0] negCond5_G256_newbasis0;
    wire [7:0] yxorb5_G256_newbasis0;
    wire [7:0] ny5_G256_newbasis0;
    wire [7:0] tempyIntoNegCond5_G256_newbasis0;
    wire [7:0] y5_G256_newbasis0;
    wire [7:0] x5_G256_newbasis0;
    wire [7:0] tempy6_G256_newbasis0;
    wire [7:0] cond6_G256_newbasis0;
    wire [7:0] negCond6_G256_newbasis0;
    wire [7:0] yxorb6_G256_newbasis0;
    wire [7:0] ny6_G256_newbasis0;
    wire [7:0] tempyIntoNegCond6_G256_newbasis0;
    wire [7:0] y6_G256_newbasis0;
    wire [7:0] x6_G256_newbasis0;
    wire [7:0] tempy7_G256_newbasis0;
    wire [7:0] cond7_G256_newbasis0;
    wire [7:0] negCond7_G256_newbasis0;
    wire [7:0] yxorb7_G256_newbasis0;
    wire [7:0] ny7_G256_newbasis0;
    wire [7:0] tempyIntoNegCond7_G256_newbasis0;
    wire [7:0] y7_G256_newbasis0;
    wire [7:0] x7_G256_newbasis0;
    wire [7:0] tempy8_G256_newbasis0;
    wire [7:0] cond8_G256_newbasis0;
    wire [7:0] negCond8_G256_newbasis0;
    wire [7:0] yxorb8_G256_newbasis0;
    wire [7:0] ny8_G256_newbasis0;
    wire [7:0] tempyIntoNegCond8_G256_newbasis0;
    wire [7:0] y8_G256_newbasis0;
    wire [7:0] x8_G256_newbasis0;
    wire [7:0] t2;
    wire [7:0] a0_0_G256_inv0;
    wire [7:0] a0_G256_inv0;
    wire [7:0] b0_G256_inv0;
    wire [7:0] a0xorb0_G256_inv0;
    wire [7:0] a0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls2_G16_sq_scl0_G256_inv0;
    wire [7:0] c0_G256_inv0;
    wire [7:0] a0_0_G16_mul0_G256_inv0;
    wire [7:0] a0_G16_mul0_G256_inv0;
    wire [7:0] b0_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G16_mul0_G256_inv0;
    wire [7:0] c0_G16_mul0_G256_inv0;
    wire [7:0] d0_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] e0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] e0_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] e01_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] e0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G16_mul0_G256_inv0;
    wire [7:0] p0_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] e0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G16_mul0_G256_inv0;
    wire [7:0] q0_G16_mul0_G256_inv0;
    wire [7:0] p0ls2_G16_mul0_G256_inv0;
    wire [7:0] d0_G256_inv0;
    wire [7:0] c0xord0_G256_inv0;
    wire [7:0] a0_0_G16_inv0_G256_inv0;
    wire [7:0] a0_G16_inv0_G256_inv0;
    wire [7:0] b0_G16_inv0_G256_inv0;
    wire [7:0] a0xorb0_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] b0ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] c0_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] c0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] d0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] e0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] d0_G16_inv0_G256_inv0;
    wire [7:0] c0xord0_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] b0ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] e0_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] c0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] d0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] e0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] c0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] d0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] e0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G16_inv0_G256_inv0;
    wire [7:0] p0ls2_G16_inv0_G256_inv0;
    wire [7:0] e0_G256_inv0;
    wire [7:0] a0_0_G16_mul1_G256_inv0;
    wire [7:0] a0_G16_mul1_G256_inv0;
    wire [7:0] b0_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G16_mul1_G256_inv0;
    wire [7:0] c0_G16_mul1_G256_inv0;
    wire [7:0] d0_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] e0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] e0_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] e01_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] e0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G16_mul1_G256_inv0;
    wire [7:0] p0_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] e0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G16_mul1_G256_inv0;
    wire [7:0] q0_G16_mul1_G256_inv0;
    wire [7:0] p0ls2_G16_mul1_G256_inv0;
    wire [7:0] p0_G256_inv0;
    wire [7:0] a0_0_G16_mul2_G256_inv0;
    wire [7:0] a0_G16_mul2_G256_inv0;
    wire [7:0] b0_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G16_mul2_G256_inv0;
    wire [7:0] c0_G16_mul2_G256_inv0;
    wire [7:0] d0_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] e0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] e0_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] e01_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] e0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G16_mul2_G256_inv0;
    wire [7:0] p0_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] e0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G16_mul2_G256_inv0;
    wire [7:0] q0_G16_mul2_G256_inv0;
    wire [7:0] p0ls2_G16_mul2_G256_inv0;
    wire [7:0] q0_G256_inv0;
    wire [7:0] p0ls4_G256_inv0;
    wire [7:0] t4;
    wire [7:0] y_G256_newbasis1;
    wire [7:0] tempy1_G256_newbasis1;
    wire [7:0] cond1_G256_newbasis1;
    wire [7:0] negCond1_G256_newbasis1;
    wire [7:0] yxorb1_G256_newbasis1;
    wire [7:0] ny1_G256_newbasis1;
    wire [7:0] tempyIntoNegCond1_G256_newbasis1;
    wire [7:0] y1_G256_newbasis1;
    wire [7:0] x1_G256_newbasis1;
    wire [7:0] tempy2_G256_newbasis1;
    wire [7:0] cond2_G256_newbasis1;
    wire [7:0] negCond2_G256_newbasis1;
    wire [7:0] yxorb2_G256_newbasis1;
    wire [7:0] ny2_G256_newbasis1;
    wire [7:0] tempyIntoNegCond2_G256_newbasis1;
    wire [7:0] y2_G256_newbasis1;
    wire [7:0] x2_G256_newbasis1;
    wire [7:0] tempy3_G256_newbasis1;
    wire [7:0] cond3_G256_newbasis1;
    wire [7:0] negCond3_G256_newbasis1;
    wire [7:0] yxorb3_G256_newbasis1;
    wire [7:0] ny3_G256_newbasis1;
    wire [7:0] tempyIntoNegCond3_G256_newbasis1;
    wire [7:0] y3_G256_newbasis1;
    wire [7:0] x3_G256_newbasis1;
    wire [7:0] tempy4_G256_newbasis1;
    wire [7:0] cond4_G256_newbasis1;
    wire [7:0] negCond4_G256_newbasis1;
    wire [7:0] yxorb4_G256_newbasis1;
    wire [7:0] ny4_G256_newbasis1;
    wire [7:0] tempyIntoNegCond4_G256_newbasis1;
    wire [7:0] y4_G256_newbasis1;
    wire [7:0] x4_G256_newbasis1;
    wire [7:0] tempy5_G256_newbasis1;
    wire [7:0] cond5_G256_newbasis1;
    wire [7:0] negCond5_G256_newbasis1;
    wire [7:0] yxorb5_G256_newbasis1;
    wire [7:0] ny5_G256_newbasis1;
    wire [7:0] tempyIntoNegCond5_G256_newbasis1;
    wire [7:0] y5_G256_newbasis1;
    wire [7:0] x5_G256_newbasis1;
    wire [7:0] tempy6_G256_newbasis1;
    wire [7:0] cond6_G256_newbasis1;
    wire [7:0] negCond6_G256_newbasis1;
    wire [7:0] yxorb6_G256_newbasis1;
    wire [7:0] ny6_G256_newbasis1;
    wire [7:0] tempyIntoNegCond6_G256_newbasis1;
    wire [7:0] y6_G256_newbasis1;
    wire [7:0] x6_G256_newbasis1;
    wire [7:0] tempy7_G256_newbasis1;
    wire [7:0] cond7_G256_newbasis1;
    wire [7:0] negCond7_G256_newbasis1;
    wire [7:0] yxorb7_G256_newbasis1;
    wire [7:0] ny7_G256_newbasis1;
    wire [7:0] tempyIntoNegCond7_G256_newbasis1;
    wire [7:0] y7_G256_newbasis1;
    wire [7:0] x7_G256_newbasis1;
    wire [7:0] tempy8_G256_newbasis1;
    wire [7:0] cond8_G256_newbasis1;
    wire [7:0] negCond8_G256_newbasis1;
    wire [7:0] yxorb8_G256_newbasis1;
    wire [7:0] ny8_G256_newbasis1;
    wire [7:0] tempyIntoNegCond8_G256_newbasis1;
    wire [7:0] y8_G256_newbasis1;
    wire [7:0] x8_G256_newbasis1;
    wire [7:0] t6;

    assign dec_99_inp = dec_99;
    assign dec_88_inp = dec_88;
    assign dec_45_inp = dec_45;
    assign dec_158_inp = dec_158;
    assign dec_11_inp = dec_11;
    assign dec_220_inp = dec_220;
    assign dec_36_inp = dec_36;
    assign dec_3_inp = dec_3;
    assign dec_2_inp = dec_2;
    assign dec_12_inp = dec_12;
    assign dec_15_inp = dec_15;
    assign dec_4_inp = dec_4;
    assign dec_240_inp = dec_240;
    assign dec_152_inp = dec_152;
    assign dec_243_inp = dec_243;
    assign dec_242_inp = dec_242;
    assign dec_72_inp = dec_72;
    assign dec_9_inp = dec_9;
    assign dec_129_inp = dec_129;
    assign dec_169_inp = dec_169;
    assign dec_255_inp = dec_255;
    assign dec_1_inp = dec_1;
    assign dec_0_inp = dec_0;
    assign t_inp = t;
    assign y_G256_newbasis0 = dec_0_inp;
    assign tempy1_G256_newbasis0 = y_G256_newbasis0;
    assign cond1_G256_newbasis0 = (t_inp & dec_1_inp);
    assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
    assign yxorb1_G256_newbasis0 = (y_G256_newbasis0 ^ dec_255_inp);
    assign ny1_G256_newbasis0 = (cond1_G256_newbasis0 * yxorb1_G256_newbasis0);
    assign tempyIntoNegCond1_G256_newbasis0 = (tempy1_G256_newbasis0 * negCond1_G256_newbasis0);
    assign y1_G256_newbasis0 = (ny1_G256_newbasis0 + tempyIntoNegCond1_G256_newbasis0);
    assign x1_G256_newbasis0 = (t_inp >> dec_1_inp);
    assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
    assign cond2_G256_newbasis0 = (x1_G256_newbasis0 & dec_1_inp);
    assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
    assign yxorb2_G256_newbasis0 = (y1_G256_newbasis0 ^ dec_169_inp);
    assign ny2_G256_newbasis0 = (cond2_G256_newbasis0 * yxorb2_G256_newbasis0);
    assign tempyIntoNegCond2_G256_newbasis0 = (tempy2_G256_newbasis0 * negCond2_G256_newbasis0);
    assign y2_G256_newbasis0 = (ny2_G256_newbasis0 + tempyIntoNegCond2_G256_newbasis0);
    assign x2_G256_newbasis0 = (x1_G256_newbasis0 >> dec_1_inp);
    assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
    assign cond3_G256_newbasis0 = (x2_G256_newbasis0 & dec_1_inp);
    assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
    assign yxorb3_G256_newbasis0 = (y2_G256_newbasis0 ^ dec_129_inp);
    assign ny3_G256_newbasis0 = (cond3_G256_newbasis0 * yxorb3_G256_newbasis0);
    assign tempyIntoNegCond3_G256_newbasis0 = (tempy3_G256_newbasis0 * negCond3_G256_newbasis0);
    assign y3_G256_newbasis0 = (ny3_G256_newbasis0 + tempyIntoNegCond3_G256_newbasis0);
    assign x3_G256_newbasis0 = (x2_G256_newbasis0 >> dec_1_inp);
    assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
    assign cond4_G256_newbasis0 = (x3_G256_newbasis0 & dec_1_inp);
    assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
    assign yxorb4_G256_newbasis0 = (y3_G256_newbasis0 ^ dec_9_inp);
    assign ny4_G256_newbasis0 = (cond4_G256_newbasis0 * yxorb4_G256_newbasis0);
    assign tempyIntoNegCond4_G256_newbasis0 = (tempy4_G256_newbasis0 * negCond4_G256_newbasis0);
    assign y4_G256_newbasis0 = (ny4_G256_newbasis0 + tempyIntoNegCond4_G256_newbasis0);
    assign x4_G256_newbasis0 = (x3_G256_newbasis0 >> dec_1_inp);
    assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
    assign cond5_G256_newbasis0 = (x4_G256_newbasis0 & dec_1_inp);
    assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
    assign yxorb5_G256_newbasis0 = (y4_G256_newbasis0 ^ dec_72_inp);
    assign ny5_G256_newbasis0 = (cond5_G256_newbasis0 * yxorb5_G256_newbasis0);
    assign tempyIntoNegCond5_G256_newbasis0 = (tempy5_G256_newbasis0 * negCond5_G256_newbasis0);
    assign y5_G256_newbasis0 = (ny5_G256_newbasis0 + tempyIntoNegCond5_G256_newbasis0);
    assign x5_G256_newbasis0 = (x4_G256_newbasis0 >> dec_1_inp);
    assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
    assign cond6_G256_newbasis0 = (x5_G256_newbasis0 & dec_1_inp);
    assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
    assign yxorb6_G256_newbasis0 = (y5_G256_newbasis0 ^ dec_242_inp);
    assign ny6_G256_newbasis0 = (cond6_G256_newbasis0 * yxorb6_G256_newbasis0);
    assign tempyIntoNegCond6_G256_newbasis0 = (tempy6_G256_newbasis0 * negCond6_G256_newbasis0);
    assign y6_G256_newbasis0 = (ny6_G256_newbasis0 + tempyIntoNegCond6_G256_newbasis0);
    assign x6_G256_newbasis0 = (x5_G256_newbasis0 >> dec_1_inp);
    assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
    assign cond7_G256_newbasis0 = (x6_G256_newbasis0 & dec_1_inp);
    assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
    assign yxorb7_G256_newbasis0 = (y6_G256_newbasis0 ^ dec_243_inp);
    assign ny7_G256_newbasis0 = (cond7_G256_newbasis0 * yxorb7_G256_newbasis0);
    assign tempyIntoNegCond7_G256_newbasis0 = (tempy7_G256_newbasis0 * negCond7_G256_newbasis0);
    assign y7_G256_newbasis0 = (ny7_G256_newbasis0 + tempyIntoNegCond7_G256_newbasis0);
    assign x7_G256_newbasis0 = (x6_G256_newbasis0 >> dec_1_inp);
    assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
    assign cond8_G256_newbasis0 = (x7_G256_newbasis0 & dec_1_inp);
    assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
    assign yxorb8_G256_newbasis0 = (y7_G256_newbasis0 ^ dec_152_inp);
    assign ny8_G256_newbasis0 = (cond8_G256_newbasis0 * yxorb8_G256_newbasis0);
    assign tempyIntoNegCond8_G256_newbasis0 = (tempy8_G256_newbasis0 * negCond8_G256_newbasis0);
    assign y8_G256_newbasis0 = (ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0);
    assign x8_G256_newbasis0 = (x7_G256_newbasis0 >> dec_1_inp);
    assign t2 = y8_G256_newbasis0;
    assign a0_0_G256_inv0 = (t2 & dec_240_inp);
    assign a0_G256_inv0 = (a0_0_G256_inv0 >> dec_4_inp);
    assign b0_G256_inv0 = (t2 & dec_15_inp);
    assign a0xorb0_G256_inv0 = (a0_G256_inv0 ^ b0_G256_inv0);
    assign a0_0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_12_inp);
    assign a0_G16_sq_scl0_G256_inv0 = (a0_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign b0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_3_inp);
    assign p0_0_G16_sq_scl0_G256_inv0 = (a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b0_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_G16_sq_scl0_G256_inv0 = (p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p0ls2_G16_sq_scl0_G256_inv0 = (p0_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign c0_G256_inv0 = (p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0);
    assign a0_0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign a0_G16_mul0_G256_inv0 = (a0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c0_G16_mul0_G256_inv0 = (c0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0);
    assign cxord_0_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0);
    assign a0_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul0_G256_inv0 = (a0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul0_G256_inv0 = (c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ d0_G4_mul0_G16_mul0_G256_inv0);
    assign e0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0 & cxord_0_G4_mul0_G16_mul0_G256_inv0);
    assign p0_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 & c0_G4_mul0_G16_mul0_G256_inv0);
    assign p0_G4_mul0_G16_mul0_G256_inv0 = (p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign q0_0_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0 & d0_G4_mul0_G16_mul0_G256_inv0);
    assign q0_G4_mul0_G16_mul0_G256_inv0 = (q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = (p0_G4_mul0_G16_mul0_G256_inv0 << dec_1_inp);
    assign e0_G16_mul0_G256_inv0 = (p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
    assign q0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0);
    assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p0_G4_scl_N0_G16_mul0_G256_inv0 << dec_1_inp);
    assign e01_G16_mul0_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0);
    assign a0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul0_G256_inv0 = (a0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul0_G256_inv0 = (c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ b0_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ d0_G4_mul1_G16_mul0_G256_inv0);
    assign e0_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0 & cxord_0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 & c0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G4_mul1_G16_mul0_G256_inv0 = (p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign q0_0_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0 & d0_G4_mul1_G16_mul0_G256_inv0);
    assign q0_G4_mul1_G16_mul0_G256_inv0 = (q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = (p0_G4_mul1_G16_mul0_G256_inv0 << dec_1_inp);
    assign p0_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G16_mul0_G256_inv0 = (p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign a0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul0_G256_inv0 = (a0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul0_G256_inv0 = (c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ b0_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ d0_G4_mul2_G16_mul0_G256_inv0);
    assign e0_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0 & cxord_0_G4_mul2_G16_mul0_G256_inv0);
    assign p0_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 & c0_G4_mul2_G16_mul0_G256_inv0);
    assign p0_G4_mul2_G16_mul0_G256_inv0 = (p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0 & d0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G4_mul2_G16_mul0_G256_inv0 = (q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = (p0_G4_mul2_G16_mul0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G16_mul0_G256_inv0 = (q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign p0ls2_G16_mul0_G256_inv0 = (p0_G16_mul0_G256_inv0 << dec_2_inp);
    assign d0_G256_inv0 = (p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0);
    assign c0xord0_G256_inv0 = (c0_G256_inv0 ^ d0_G256_inv0);
    assign a0_0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_12_inp);
    assign a0_G16_inv0_G256_inv0 = (a0_0_G16_inv0_G256_inv0 >> dec_2_inp);
    assign b0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_3_inp);
    assign a0xorb0_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 ^ b0_G16_inv0_G256_inv0);
    assign a0_0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq2_G16_inv0_G256_inv0 = (a0_0_G4_sq2_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = (b0_G4_sq2_G16_inv0_G256_inv0 << dec_1_inp);
    assign c0_0_G16_inv0_G256_inv0 = (b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0);
    assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
    assign q0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0);
    assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p0_G4_scl_N1_G16_inv0_G256_inv0 << dec_1_inp);
    assign c0_G16_inv0_G256_inv0 = (p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0);
    assign a0_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul3_G16_inv0_G256_inv0 = (a0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul3_G16_inv0_G256_inv0 = (c0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ b0_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ d0_G4_mul3_G16_inv0_G256_inv0);
    assign e0_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0 & cxord_0_G4_mul3_G16_inv0_G256_inv0);
    assign p0_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 & c0_G4_mul3_G16_inv0_G256_inv0);
    assign p0_G4_mul3_G16_inv0_G256_inv0 = (p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign q0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0 & d0_G4_mul3_G16_inv0_G256_inv0);
    assign q0_G4_mul3_G16_inv0_G256_inv0 = (q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = (p0_G4_mul3_G16_inv0_G256_inv0 << dec_1_inp);
    assign d0_G16_inv0_G256_inv0 = (p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0);
    assign c0xord0_G16_inv0_G256_inv0 = (c0_G16_inv0_G256_inv0 ^ d0_G16_inv0_G256_inv0);
    assign a0_0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq3_G16_inv0_G256_inv0 = (a0_0_G4_sq3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = (b0_G4_sq3_G16_inv0_G256_inv0 << dec_1_inp);
    assign e0_G16_inv0_G256_inv0 = (b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0);
    assign a0_0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul4_G16_inv0_G256_inv0 = (a0_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul4_G16_inv0_G256_inv0 = (c0_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ d0_G4_mul4_G16_inv0_G256_inv0);
    assign e0_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & cxord_0_G4_mul4_G16_inv0_G256_inv0);
    assign p0_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & c0_G4_mul4_G16_inv0_G256_inv0);
    assign p0_G4_mul4_G16_inv0_G256_inv0 = (p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign q0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & d0_G4_mul4_G16_inv0_G256_inv0);
    assign q0_G4_mul4_G16_inv0_G256_inv0 = (q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = (p0_G4_mul4_G16_inv0_G256_inv0 << dec_1_inp);
    assign p0_G16_inv0_G256_inv0 = (p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0);
    assign a0_0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul5_G16_inv0_G256_inv0 = (a0_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul5_G16_inv0_G256_inv0 = (c0_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ b0_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ d0_G4_mul5_G16_inv0_G256_inv0);
    assign e0_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & cxord_0_G4_mul5_G16_inv0_G256_inv0);
    assign p0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & c0_G4_mul5_G16_inv0_G256_inv0);
    assign p0_G4_mul5_G16_inv0_G256_inv0 = (p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign q0_0_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & d0_G4_mul5_G16_inv0_G256_inv0);
    assign q0_G4_mul5_G16_inv0_G256_inv0 = (q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = (p0_G4_mul5_G16_inv0_G256_inv0 << dec_1_inp);
    assign q0_G16_inv0_G256_inv0 = (p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0);
    assign p0ls2_G16_inv0_G256_inv0 = (p0_G16_inv0_G256_inv0 << dec_2_inp);
    assign e0_G256_inv0 = (p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0);
    assign a0_0_G16_mul1_G256_inv0 = (e0_G256_inv0 & dec_12_inp);
    assign a0_G16_mul1_G256_inv0 = (a0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul1_G256_inv0 = (e0_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c0_G16_mul1_G256_inv0 = (c0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0);
    assign cxord_0_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0);
    assign a0_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul1_G256_inv0 = (a0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul1_G256_inv0 = (c0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ b0_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ d0_G4_mul0_G16_mul1_G256_inv0);
    assign e0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & cxord_0_G4_mul0_G16_mul1_G256_inv0);
    assign p0_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & c0_G4_mul0_G16_mul1_G256_inv0);
    assign p0_G4_mul0_G16_mul1_G256_inv0 = (p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign q0_0_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & d0_G4_mul0_G16_mul1_G256_inv0);
    assign q0_G4_mul0_G16_mul1_G256_inv0 = (q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = (p0_G4_mul0_G16_mul1_G256_inv0 << dec_1_inp);
    assign e0_G16_mul1_G256_inv0 = (p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
    assign q0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0);
    assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p0_G4_scl_N0_G16_mul1_G256_inv0 << dec_1_inp);
    assign e01_G16_mul1_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0);
    assign a0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul1_G256_inv0 = (a0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul1_G256_inv0 = (c0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ b0_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ d0_G4_mul1_G16_mul1_G256_inv0);
    assign e0_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & cxord_0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & c0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G4_mul1_G16_mul1_G256_inv0 = (p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign q0_0_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & d0_G4_mul1_G16_mul1_G256_inv0);
    assign q0_G4_mul1_G16_mul1_G256_inv0 = (q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = (p0_G4_mul1_G16_mul1_G256_inv0 << dec_1_inp);
    assign p0_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G16_mul1_G256_inv0 = (p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign a0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul1_G256_inv0 = (a0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul1_G256_inv0 = (c0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ d0_G4_mul2_G16_mul1_G256_inv0);
    assign e0_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & cxord_0_G4_mul2_G16_mul1_G256_inv0);
    assign p0_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & c0_G4_mul2_G16_mul1_G256_inv0);
    assign p0_G4_mul2_G16_mul1_G256_inv0 = (p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & d0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G4_mul2_G16_mul1_G256_inv0 = (q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = (p0_G4_mul2_G16_mul1_G256_inv0 << dec_1_inp);
    assign q0_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G16_mul1_G256_inv0 = (q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign p0ls2_G16_mul1_G256_inv0 = (p0_G16_mul1_G256_inv0 << dec_2_inp);
    assign p0_G256_inv0 = (p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0);
    assign a0_0_G16_mul2_G256_inv0 = (e0_G256_inv0 & dec_12_inp);
    assign a0_G16_mul2_G256_inv0 = (a0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul2_G256_inv0 = (e0_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign c0_G16_mul2_G256_inv0 = (c0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0);
    assign cxord_0_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0);
    assign a0_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul2_G256_inv0 = (a0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul2_G256_inv0 = (c0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ d0_G4_mul0_G16_mul2_G256_inv0);
    assign e0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & cxord_0_G4_mul0_G16_mul2_G256_inv0);
    assign p0_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & c0_G4_mul0_G16_mul2_G256_inv0);
    assign p0_G4_mul0_G16_mul2_G256_inv0 = (p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign q0_0_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & d0_G4_mul0_G16_mul2_G256_inv0);
    assign q0_G4_mul0_G16_mul2_G256_inv0 = (q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = (p0_G4_mul0_G16_mul2_G256_inv0 << dec_1_inp);
    assign e0_G16_mul2_G256_inv0 = (p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
    assign q0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0);
    assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p0_G4_scl_N0_G16_mul2_G256_inv0 << dec_1_inp);
    assign e01_G16_mul2_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0);
    assign a0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul2_G256_inv0 = (a0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul2_G256_inv0 = (c0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ d0_G4_mul1_G16_mul2_G256_inv0);
    assign e0_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & cxord_0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & c0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G4_mul1_G16_mul2_G256_inv0 = (p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign q0_0_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & d0_G4_mul1_G16_mul2_G256_inv0);
    assign q0_G4_mul1_G16_mul2_G256_inv0 = (q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = (p0_G4_mul1_G16_mul2_G256_inv0 << dec_1_inp);
    assign p0_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G16_mul2_G256_inv0 = (p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign a0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul2_G256_inv0 = (a0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul2_G256_inv0 = (c0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ d0_G4_mul2_G16_mul2_G256_inv0);
    assign e0_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & cxord_0_G4_mul2_G16_mul2_G256_inv0);
    assign p0_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & c0_G4_mul2_G16_mul2_G256_inv0);
    assign p0_G4_mul2_G16_mul2_G256_inv0 = (p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & d0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G4_mul2_G16_mul2_G256_inv0 = (q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = (p0_G4_mul2_G16_mul2_G256_inv0 << dec_1_inp);
    assign q0_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G16_mul2_G256_inv0 = (q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign p0ls2_G16_mul2_G256_inv0 = (p0_G16_mul2_G256_inv0 << dec_2_inp);
    assign q0_G256_inv0 = (p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0);
    assign p0ls4_G256_inv0 = (p0_G256_inv0 << dec_4_inp);
    assign t4 = (p0ls4_G256_inv0 | q0_G256_inv0);
    assign y_G256_newbasis1 = dec_0_inp;
    assign tempy1_G256_newbasis1 = y_G256_newbasis1;
    assign cond1_G256_newbasis1 = (t4 & dec_1_inp);
    assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
    assign yxorb1_G256_newbasis1 = (y_G256_newbasis1 ^ dec_36_inp);
    assign ny1_G256_newbasis1 = (cond1_G256_newbasis1 * yxorb1_G256_newbasis1);
    assign tempyIntoNegCond1_G256_newbasis1 = (tempy1_G256_newbasis1 * negCond1_G256_newbasis1);
    assign y1_G256_newbasis1 = (ny1_G256_newbasis1 + tempyIntoNegCond1_G256_newbasis1);
    assign x1_G256_newbasis1 = (t4 >> dec_1_inp);
    assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
    assign cond2_G256_newbasis1 = (x1_G256_newbasis1 & dec_1_inp);
    assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
    assign yxorb2_G256_newbasis1 = (y1_G256_newbasis1 ^ dec_3_inp);
    assign ny2_G256_newbasis1 = (cond2_G256_newbasis1 * yxorb2_G256_newbasis1);
    assign tempyIntoNegCond2_G256_newbasis1 = (tempy2_G256_newbasis1 * negCond2_G256_newbasis1);
    assign y2_G256_newbasis1 = (ny2_G256_newbasis1 + tempyIntoNegCond2_G256_newbasis1);
    assign x2_G256_newbasis1 = (x1_G256_newbasis1 >> dec_1_inp);
    assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
    assign cond3_G256_newbasis1 = (x2_G256_newbasis1 & dec_1_inp);
    assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
    assign yxorb3_G256_newbasis1 = (y2_G256_newbasis1 ^ dec_4_inp);
    assign ny3_G256_newbasis1 = (cond3_G256_newbasis1 * yxorb3_G256_newbasis1);
    assign tempyIntoNegCond3_G256_newbasis1 = (tempy3_G256_newbasis1 * negCond3_G256_newbasis1);
    assign y3_G256_newbasis1 = (ny3_G256_newbasis1 + tempyIntoNegCond3_G256_newbasis1);
    assign x3_G256_newbasis1 = (x2_G256_newbasis1 >> dec_1_inp);
    assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
    assign cond4_G256_newbasis1 = (x3_G256_newbasis1 & dec_1_inp);
    assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
    assign yxorb4_G256_newbasis1 = (y3_G256_newbasis1 ^ dec_220_inp);
    assign ny4_G256_newbasis1 = (cond4_G256_newbasis1 * yxorb4_G256_newbasis1);
    assign tempyIntoNegCond4_G256_newbasis1 = (tempy4_G256_newbasis1 * negCond4_G256_newbasis1);
    assign y4_G256_newbasis1 = (ny4_G256_newbasis1 + tempyIntoNegCond4_G256_newbasis1);
    assign x4_G256_newbasis1 = (x3_G256_newbasis1 >> dec_1_inp);
    assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
    assign cond5_G256_newbasis1 = (x4_G256_newbasis1 & dec_1_inp);
    assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
    assign yxorb5_G256_newbasis1 = (y4_G256_newbasis1 ^ dec_11_inp);
    assign ny5_G256_newbasis1 = (cond5_G256_newbasis1 * yxorb5_G256_newbasis1);
    assign tempyIntoNegCond5_G256_newbasis1 = (tempy5_G256_newbasis1 * negCond5_G256_newbasis1);
    assign y5_G256_newbasis1 = (ny5_G256_newbasis1 + tempyIntoNegCond5_G256_newbasis1);
    assign x5_G256_newbasis1 = (x4_G256_newbasis1 >> dec_1_inp);
    assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
    assign cond6_G256_newbasis1 = (x5_G256_newbasis1 & dec_1_inp);
    assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
    assign yxorb6_G256_newbasis1 = (y5_G256_newbasis1 ^ dec_158_inp);
    assign ny6_G256_newbasis1 = (cond6_G256_newbasis1 * yxorb6_G256_newbasis1);
    assign tempyIntoNegCond6_G256_newbasis1 = (tempy6_G256_newbasis1 * negCond6_G256_newbasis1);
    assign y6_G256_newbasis1 = (ny6_G256_newbasis1 + tempyIntoNegCond6_G256_newbasis1);
    assign x6_G256_newbasis1 = (x5_G256_newbasis1 >> dec_1_inp);
    assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
    assign cond7_G256_newbasis1 = (x6_G256_newbasis1 & dec_1_inp);
    assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
    assign yxorb7_G256_newbasis1 = (y6_G256_newbasis1 ^ dec_45_inp);
    assign ny7_G256_newbasis1 = (cond7_G256_newbasis1 * yxorb7_G256_newbasis1);
    assign tempyIntoNegCond7_G256_newbasis1 = (tempy7_G256_newbasis1 * negCond7_G256_newbasis1);
    assign y7_G256_newbasis1 = (ny7_G256_newbasis1 + tempyIntoNegCond7_G256_newbasis1);
    assign x7_G256_newbasis1 = (x6_G256_newbasis1 >> dec_1_inp);
    assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
    assign cond8_G256_newbasis1 = (x7_G256_newbasis1 & dec_1_inp);
    assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
    assign yxorb8_G256_newbasis1 = (y7_G256_newbasis1 ^ dec_88_inp);
    assign ny8_G256_newbasis1 = (cond8_G256_newbasis1 * yxorb8_G256_newbasis1);
    assign tempyIntoNegCond8_G256_newbasis1 = (tempy8_G256_newbasis1 * negCond8_G256_newbasis1);
    assign y8_G256_newbasis1 = (ny8_G256_newbasis1 + tempyIntoNegCond8_G256_newbasis1);
    assign x8_G256_newbasis1 = (x7_G256_newbasis1 >> dec_1_inp);
    assign t6 = y8_G256_newbasis1;

    always @(posedge clk) begin
        y <= (t6 ^ dec_99_inp);
    end

endmodule

