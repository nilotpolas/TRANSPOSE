`timescale 1 ns / 1 ps


module aes_main_AddRoundKey_InversMixColumn
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  n,
  word_address0,
  word_ce0,
  word_q0,
  word_address1,
  word_ce1,
  word_q1,
  statemt_address0,
  statemt_ce0,
  statemt_we0,
  statemt_d0,
  statemt_q0,
  statemt_address1,
  statemt_ce1,
  statemt_we1,
  statemt_d1,
  statemt_q1
);

  parameter ap_ST_fsm_state1 = 12'd1;
  parameter ap_ST_fsm_state2 = 12'd2;
  parameter ap_ST_fsm_state3 = 12'd4;
  parameter ap_ST_fsm_state4 = 12'd8;
  parameter ap_ST_fsm_state5 = 12'd16;
  parameter ap_ST_fsm_state6 = 12'd32;
  parameter ap_ST_fsm_state7 = 12'd64;
  parameter ap_ST_fsm_state8 = 12'd128;
  parameter ap_ST_fsm_state9 = 12'd256;
  parameter ap_ST_fsm_state10 = 12'd512;
  parameter ap_ST_fsm_state11 = 12'd1024;
  parameter ap_ST_fsm_state12 = 12'd2048;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  input [3:0] n;
  output [8:0] word_address0;
  output word_ce0;
  input [31:0] word_q0;
  output [8:0] word_address1;
  output word_ce1;
  input [31:0] word_q1;
  output [4:0] statemt_address0;
  output statemt_ce0;
  output statemt_we0;
  output [31:0] statemt_d0;
  input [31:0] statemt_q0;
  output [4:0] statemt_address1;
  output statemt_ce1;
  output statemt_we1;
  output [31:0] statemt_d1;
  input [31:0] statemt_q1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [8:0] word_address0;
  reg word_ce0;
  reg [8:0] word_address1;
  reg word_ce1;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  (* fsm_encoding = "none" *)
  reg [11:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [31:0] grp_fu_309_p2;
  reg [31:0] reg_341;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state4;
  wire [31:0] grp_fu_315_p2;
  reg [31:0] reg_346;
  wire [5:0] mul_fu_351_p3;
  reg [5:0] mul_reg_1299;
  wire [5:0] add_ln514_fu_383_p2;
  reg [5:0] add_ln514_reg_1307;
  wire ap_CS_fsm_state2;
  wire [0:0] icmp_ln510_fu_371_p2;
  wire [3:0] shl_ln_fu_412_p3;
  reg [3:0] shl_ln_reg_1322;
  reg [4:0] statemt_addr_reg_1328;
  reg [4:0] statemt_addr_12_reg_1333;
  reg [4:0] statemt_addr_13_reg_1355;
  reg [4:0] statemt_addr_14_reg_1360;
  wire [2:0] add_ln519_fu_500_p2;
  reg [2:0] add_ln519_reg_1368;
  wire ap_CS_fsm_state6;
  wire [1:0] empty_86_fu_506_p1;
  reg [1:0] empty_86_reg_1373;
  wire [0:0] icmp_ln519_fu_494_p2;
  wire [3:0] tmp_s_fu_510_p3;
  reg [3:0] tmp_s_reg_1379;
  wire [4:0] zext_ln520_fu_518_p1;
  reg [4:0] zext_ln520_reg_1384;
  wire [2:0] add_ln459_fu_537_p2;
  reg [2:0] add_ln459_reg_1399;
  wire ap_CS_fsm_state7;
  wire [63:0] zext_ln446_fu_548_p1;
  reg [63:0] zext_ln446_reg_1404;
  wire [0:0] icmp_ln520_fu_531_p2;
  wire [1:0] trunc_ln459_fu_553_p1;
  reg [1:0] trunc_ln459_reg_1414;
  reg [31:0] statemt_load_29_reg_1425;
  wire ap_CS_fsm_state8;
  wire [31:0] xor_ln528_3_fu_919_p2;
  reg [31:0] xor_ln528_3_reg_1440;
  wire [3:0] shl_ln1_fu_1243_p3;
  reg [3:0] shl_ln1_reg_1448;
  wire ap_CS_fsm_state10;
  wire [0:0] icmp_ln531_fu_1227_p2;
  wire [63:0] zext_ln535_fu_1251_p1;
  reg [63:0] zext_ln535_reg_1454;
  wire [63:0] zext_ln536_fu_1262_p1;
  reg [63:0] zext_ln536_reg_1464;
  wire [63:0] zext_ln537_fu_1277_p1;
  reg [63:0] zext_ln537_reg_1474;
  wire ap_CS_fsm_state11;
  wire [63:0] zext_ln538_fu_1287_p1;
  reg [63:0] zext_ln538_reg_1484;
  reg [4:0] ret_address0;
  reg ret_ce0;
  reg ret_we0;
  wire [31:0] ret_d0;
  wire [31:0] ret_q0;
  reg [4:0] ret_address1;
  reg ret_ce1;
  wire [31:0] ret_q1;
  reg [2:0] i_6_reg_298;
  wire ap_CS_fsm_state9;
  wire [63:0] zext_ln514_fu_388_p1;
  wire [63:0] zext_ln515_1_fu_403_p1;
  wire [63:0] zext_ln514_1_fu_420_p1;
  wire [63:0] zext_ln515_fu_431_p1;
  wire [63:0] zext_ln516_1_fu_455_p1;
  wire [63:0] zext_ln517_1_fu_466_p1;
  wire [63:0] zext_ln516_fu_476_p1;
  wire [63:0] zext_ln517_fu_486_p1;
  wire [63:0] zext_ln459_fu_590_p1;
  wire [63:0] zext_ln475_fu_897_p1;
  wire [63:0] zext_ln488_fu_914_p1;
  wire ap_CS_fsm_state12;
  reg [2:0] j_fu_82;
  wire [2:0] add_ln510_fu_377_p2;
  reg [2:0] j_4_fu_90;
  reg [2:0] i_fu_94;
  wire [2:0] add_ln531_fu_1233_p2;
  wire ap_CS_fsm_state5;
  wire [5:0] zext_ln510_fu_367_p1;
  wire [7:0] zext_ln514_3_fu_393_p1;
  wire [7:0] add_ln515_fu_397_p2;
  wire [1:0] trunc_ln514_fu_408_p1;
  wire [3:0] or_ln515_fu_425_p2;
  wire [8:0] zext_ln514_2_fu_446_p1;
  wire [8:0] add_ln516_fu_449_p2;
  wire [8:0] add_ln517_fu_460_p2;
  wire [3:0] or_ln516_fu_471_p2;
  wire [3:0] or_ln517_fu_481_p2;
  wire [3:0] zext_ln520_1_fu_527_p1;
  wire [3:0] add_ln446_fu_543_p2;
  wire [2:0] zext_ln459_1_fu_557_p1;
  wire [0:0] empty_88_fu_561_p2;
  wire [2:0] empty_89_fu_567_p2;
  wire [2:0] iv_rem_fu_573_p3;
  wire [4:0] zext_ln459_2_fu_581_p1;
  wire [4:0] add_ln459_1_fu_585_p2;
  wire [23:0] grp_fu_321_p4;
  wire [31:0] and_ln_fu_599_p3;
  wire [29:0] trunc_ln448_fu_613_p1;
  wire [30:0] trunc_ln_fu_617_p3;
  wire [0:0] icmp_ln447_fu_607_p2;
  wire [30:0] xor_ln447_fu_625_p2;
  wire [30:0] select_ln447_fu_631_p3;
  wire [30:0] trunc_ln449_fu_639_p1;
  wire [30:0] xor_ln450_fu_643_p2;
  wire [23:0] tmp_21_fu_649_p4;
  wire [31:0] and_ln1_fu_659_p3;
  wire [30:0] shl_ln452_fu_673_p2;
  wire [0:0] icmp_ln451_fu_667_p2;
  wire [30:0] xor_ln451_fu_679_p2;
  wire [30:0] select_ln451_fu_685_p3;
  wire [30:0] xor_ln454_fu_693_p2;
  wire [23:0] tmp_22_fu_707_p4;
  wire [31:0] and_ln2_fu_717_p3;
  wire [31:0] x_assign_2_fu_699_p3;
  wire [0:0] icmp_ln455_fu_725_p2;
  wire [31:0] xor_ln456_fu_731_p2;
  wire [29:0] trunc_ln445_fu_745_p1;
  wire [23:0] grp_fu_331_p4;
  wire [31:0] and_ln3_fu_757_p3;
  wire [30:0] trunc_ln1_fu_749_p3;
  wire [0:0] icmp_ln460_fu_765_p2;
  wire [30:0] xor_ln461_fu_771_p2;
  wire [30:0] select_ln460_fu_777_p3;
  wire [23:0] tmp_24_fu_785_p4;
  wire [31:0] and_ln4_fu_795_p3;
  wire [30:0] shl_ln464_fu_809_p2;
  wire [0:0] icmp_ln463_fu_803_p2;
  wire [30:0] xor_ln463_fu_815_p2;
  wire [30:0] select_ln463_fu_821_p3;
  wire [30:0] trunc_ln465_fu_829_p1;
  wire [30:0] xor_ln466_fu_833_p2;
  wire [23:0] tmp_25_fu_847_p4;
  wire [31:0] and_ln5_fu_857_p3;
  wire [31:0] x_assign_8_fu_839_p3;
  wire [0:0] icmp_ln467_fu_865_p2;
  wire [31:0] xor_ln468_fu_871_p2;
  wire [1:0] xor_ln475_fu_885_p2;
  wire [3:0] or_ln_fu_890_p3;
  wire [1:0] add_ln488_fu_902_p2;
  wire [3:0] or_ln1_fu_907_p3;
  wire [31:0] select_ln455_fu_737_p3;
  wire [31:0] select_ln467_fu_877_p3;
  wire [31:0] and_ln6_fu_925_p3;
  wire [29:0] trunc_ln477_fu_939_p1;
  wire [30:0] trunc_ln2_fu_943_p3;
  wire [0:0] icmp_ln476_fu_933_p2;
  wire [30:0] xor_ln476_fu_951_p2;
  wire [30:0] select_ln476_fu_957_p3;
  wire [30:0] trunc_ln478_fu_965_p1;
  wire [30:0] xor_ln479_fu_969_p2;
  wire [23:0] tmp_27_fu_981_p4;
  wire [31:0] and_ln7_fu_991_p3;
  wire [30:0] shl_ln474_fu_975_p2;
  wire [0:0] icmp_ln480_fu_999_p2;
  wire [30:0] xor_ln481_fu_1005_p2;
  wire [30:0] select_ln480_fu_1011_p3;
  wire [23:0] tmp_28_fu_1027_p4;
  wire [31:0] and_ln8_fu_1037_p3;
  wire [31:0] x_assign_s_fu_1019_p3;
  wire [0:0] icmp_ln483_fu_1045_p2;
  wire [31:0] xor_ln484_fu_1051_p2;
  wire [29:0] trunc_ln474_fu_1065_p1;
  wire [31:0] and_ln9_fu_1077_p3;
  wire [30:0] trunc_ln474_1_fu_1069_p3;
  wire [0:0] icmp_ln489_fu_1085_p2;
  wire [30:0] xor_ln490_fu_1091_p2;
  wire [30:0] select_ln489_fu_1097_p3;
  wire [23:0] tmp_30_fu_1111_p4;
  wire [31:0] and_ln10_fu_1121_p3;
  wire [30:0] shl_ln474_1_fu_1105_p2;
  wire [0:0] icmp_ln492_fu_1129_p2;
  wire [30:0] xor_ln493_fu_1135_p2;
  wire [30:0] select_ln492_fu_1141_p3;
  wire [23:0] tmp_31_fu_1157_p4;
  wire [31:0] and_ln11_fu_1167_p3;
  wire [31:0] x_assign_1_fu_1149_p3;
  wire [0:0] icmp_ln495_fu_1175_p2;
  wire [31:0] xor_ln496_fu_1181_p2;
  wire [31:0] xor_ln528_1_fu_1195_p2;
  wire [31:0] select_ln483_fu_1057_p3;
  wire [31:0] select_ln495_fu_1187_p3;
  wire [31:0] xor_ln528_4_fu_1206_p2;
  wire [31:0] xor_ln528_5_fu_1212_p2;
  wire [31:0] xor_ln528_2_fu_1200_p2;
  wire [1:0] trunc_ln535_fu_1239_p1;
  wire [3:0] or_ln536_fu_1256_p2;
  wire [3:0] or_ln537_fu_1272_p2;
  wire [3:0] or_ln538_fu_1282_p2;
  reg [11:0] ap_NS_fsm;
  reg ap_ST_fsm_state1_blk;
  wire ap_ST_fsm_state2_blk;
  wire ap_ST_fsm_state3_blk;
  wire ap_ST_fsm_state4_blk;
  wire ap_ST_fsm_state5_blk;
  wire ap_ST_fsm_state6_blk;
  wire ap_ST_fsm_state7_blk;
  wire ap_ST_fsm_state8_blk;
  wire ap_ST_fsm_state9_blk;
  wire ap_ST_fsm_state10_blk;
  wire ap_ST_fsm_state11_blk;
  wire ap_ST_fsm_state12_blk;
  wire ap_ce_reg;

  initial begin
    #0 ap_CS_fsm = 12'd1;
  end


  aes_main_AddRoundKey_InversMixColumn_ret_RAM_AUTO_1R1W
  #(
    .DataWidth(32),
    .AddressRange(32),
    .AddressWidth(5)
  )
  ret_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(ret_address0),
    .ce0(ret_ce0),
    .we0(ret_we0),
    .d0(ret_d0),
    .q0(ret_q0),
    .address1(ret_address1),
    .ce1(ret_ce1),
    .q1(ret_q1)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state6) & (icmp_ln519_fu_494_p2 == 1'd0)) begin
      i_6_reg_298 <= 3'd0;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      i_6_reg_298 <= add_ln459_reg_1399;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state6) & (icmp_ln519_fu_494_p2 == 1'd1)) begin
      i_fu_94 <= 3'd0;
    end else if((1'b1 == ap_CS_fsm_state10) & (icmp_ln531_fu_1227_p2 == 1'd0)) begin
      i_fu_94 <= add_ln531_fu_1233_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln510_fu_371_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      j_4_fu_90 <= 3'd0;
    end else if((1'b1 == ap_CS_fsm_state7) & (icmp_ln520_fu_531_p2 == 1'd1)) begin
      j_4_fu_90 <= ~add_ln519_reg_1368;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      j_fu_82 <= 3'd0;
    end else if((icmp_ln510_fu_371_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      j_fu_82 <= add_ln510_fu_377_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      add_ln459_reg_1399 <= add_ln459_fu_537_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln510_fu_371_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      add_ln514_reg_1307 <= add_ln514_fu_383_p2;
      shl_ln_reg_1322[3:2] <= shl_ln_fu_412_p3[3:2];
      statemt_addr_12_reg_1333[3:2] <= zext_ln515_fu_431_p1[3:2];
      statemt_addr_reg_1328[3:2] <= zext_ln514_1_fu_420_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      add_ln519_reg_1368 <= add_ln519_fu_500_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state6) & (icmp_ln519_fu_494_p2 == 1'd0)) begin
      empty_86_reg_1373 <= empty_86_fu_506_p1;
      tmp_s_reg_1379[3:2] <= tmp_s_fu_510_p3[3:2];
      zext_ln520_reg_1384[3:2] <= zext_ln520_fu_518_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state1) begin
      mul_reg_1299[5:2] <= mul_fu_351_p3[5:2];
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3)) begin
      reg_341 <= grp_fu_309_p2;
      reg_346 <= grp_fu_315_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state10) & (icmp_ln531_fu_1227_p2 == 1'd0)) begin
      shl_ln1_reg_1448[3:2] <= shl_ln1_fu_1243_p3[3:2];
      zext_ln535_reg_1454[3:2] <= zext_ln535_fu_1251_p1[3:2];
      zext_ln536_reg_1464[3:2] <= zext_ln536_fu_1262_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_addr_13_reg_1355[3:2] <= ~zext_ln516_fu_476_p1[3:2];
      statemt_addr_14_reg_1360[3:2] <= zext_ln517_fu_486_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      statemt_load_29_reg_1425 <= ~statemt_q0;
      xor_ln528_3_reg_1440 <= xor_ln528_3_fu_919_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state7) & (icmp_ln520_fu_531_p2 == 1'd0)) begin
      trunc_ln459_reg_1414 <= trunc_ln459_fu_553_p1;
      zext_ln446_reg_1404[3:0] <= zext_ln446_fu_548_p1[3:0];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      zext_ln537_reg_1474[3:2] <= zext_ln537_fu_1277_p1[3:2];
      zext_ln538_reg_1484[3:2] <= zext_ln538_fu_1287_p1[3:2];
    end 
  end

  assign ap_ST_fsm_state10_blk = 1'b0;
  assign ap_ST_fsm_state11_blk = 1'b0;
  assign ap_ST_fsm_state12_blk = 1'b0;

  always @(*) begin
    if(ap_start == 1'b0) begin
      ap_ST_fsm_state1_blk = 1'b1;
    end else begin
      ap_ST_fsm_state1_blk = 1'b0;
    end
  end

  assign ap_ST_fsm_state2_blk = 1'b0;
  assign ap_ST_fsm_state3_blk = 1'b0;
  assign ap_ST_fsm_state4_blk = 1'b0;
  assign ap_ST_fsm_state5_blk = 1'b0;
  assign ap_ST_fsm_state6_blk = 1'b0;
  assign ap_ST_fsm_state7_blk = 1'b0;
  assign ap_ST_fsm_state8_blk = 1'b0;
  assign ap_ST_fsm_state9_blk = 1'b0;

  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0) | (1'b1 == ap_CS_fsm_state10) & (icmp_ln531_fu_1227_p2 == 1'd1)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state10) & (icmp_ln531_fu_1227_p2 == 1'd1)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      ret_address0 = zext_ln537_fu_1277_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      ret_address0 = zext_ln536_fu_1262_p1;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      ret_address0 = zext_ln446_reg_1404;
    end else begin
      ret_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      ret_address1 = zext_ln538_fu_1287_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      ret_address1 = zext_ln535_fu_1251_p1;
    end else begin
      ret_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10)) begin
      ret_ce0 = 1'b1;
    end else begin
      ret_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10)) begin
      ret_ce1 = 1'b1;
    end else begin
      ret_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      ret_we0 = 1'b1;
    end else begin
      ret_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address0 = zext_ln538_reg_1484;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_address0 = zext_ln536_reg_1464;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = zext_ln488_fu_914_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address0 = zext_ln459_fu_590_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address0 = statemt_addr_14_reg_1360;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address0 = statemt_addr_12_reg_1333;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = zext_ln517_fu_486_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address0 = zext_ln515_fu_431_p1;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address1 = zext_ln537_reg_1474;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_address1 = zext_ln535_reg_1454;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = zext_ln475_fu_897_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address1 = zext_ln446_fu_548_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address1 = ~statemt_addr_13_reg_1355;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address1 = ~statemt_addr_reg_1328;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address1 = zext_ln516_fu_476_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address1 = ~zext_ln514_1_fu_420_p1;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7)) begin
      statemt_ce0 = 1'b1;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7)) begin
      statemt_ce1 = 1'b1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      statemt_d0 = ret_q1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_d0 = ret_q0;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d0 = reg_346;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      statemt_d1 = ret_q0;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_d1 = ret_q1;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d1 = reg_341;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11)) begin
      statemt_we0 = 1'b1;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11)) begin
      statemt_we1 = 1'b1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address0 = zext_ln517_1_fu_466_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address0 = zext_ln515_1_fu_403_p1;
    end else begin
      word_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address1 = zext_ln516_1_fu_455_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address1 = zext_ln514_fu_388_p1;
    end else begin
      word_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce0 = 1'b1;
    end else begin
      word_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce1 = 1'b1;
    end else begin
      word_ce1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((icmp_ln510_fu_371_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state4;
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      ap_ST_fsm_state6: begin
        if((1'b1 == ap_CS_fsm_state6) & (icmp_ln519_fu_494_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end
      end
      ap_ST_fsm_state7: begin
        if((1'b1 == ap_CS_fsm_state7) & (icmp_ln520_fu_531_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state10: begin
        if((1'b1 == ap_CS_fsm_state10) & (icmp_ln531_fu_1227_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state12: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign add_ln446_fu_543_p2 = zext_ln520_1_fu_527_p1 + tmp_s_reg_1379;
  assign add_ln459_1_fu_585_p2 = zext_ln459_2_fu_581_p1 + zext_ln520_reg_1384;
  assign add_ln459_fu_537_p2 = i_6_reg_298 + 3'd1;
  assign add_ln488_fu_902_p2 = $signed(trunc_ln459_reg_1414) + $signed(2'd3);
  assign add_ln510_fu_377_p2 = j_fu_82 + 3'd1;
  assign add_ln514_fu_383_p2 = zext_ln510_fu_367_p1 + mul_reg_1299;
  assign add_ln515_fu_397_p2 = zext_ln514_3_fu_393_p1 + 8'd120;
  assign add_ln516_fu_449_p2 = zext_ln514_2_fu_446_p1 + 9'd240;
  assign add_ln517_fu_460_p2 = $signed(zext_ln514_2_fu_446_p1) + $signed(9'd360);
  assign add_ln519_fu_500_p2 = ~j_4_fu_90 + (~3'd1 + 1);
  assign add_ln531_fu_1233_p2 = i_fu_94 + 3'd1;
  assign and_ln10_fu_1121_p3 = { { tmp_30_fu_1111_p4 }, { 8'd0 } };
  assign and_ln11_fu_1167_p3 = { { tmp_31_fu_1157_p4 }, { 8'd0 } };
  assign and_ln1_fu_659_p3 = { { tmp_21_fu_649_p4 }, { 8'd0 } };
  assign and_ln2_fu_717_p3 = { { tmp_22_fu_707_p4 }, { 8'd0 } };
  assign and_ln3_fu_757_p3 = { { grp_fu_331_p4 }, { 8'd0 } };
  assign and_ln4_fu_795_p3 = { { tmp_24_fu_785_p4 }, { 8'd0 } };
  assign and_ln5_fu_857_p3 = { { tmp_25_fu_847_p4 }, { 8'd0 } };
  assign and_ln6_fu_925_p3 = { { grp_fu_321_p4 }, { 8'd0 } };
  assign and_ln7_fu_991_p3 = { { tmp_27_fu_981_p4 }, { 8'd0 } };
  assign and_ln8_fu_1037_p3 = { { tmp_28_fu_1027_p4 }, { 8'd0 } };
  assign and_ln9_fu_1077_p3 = { { grp_fu_331_p4 }, { 8'd0 } };
  assign and_ln_fu_599_p3 = { { grp_fu_321_p4 }, { 8'd0 } };
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign empty_86_fu_506_p1 = j_4_fu_90[1:0];
  assign empty_88_fu_561_p2 = (add_ln459_fu_537_p2 == 3'd4)? 1'b1 : 1'b0;
  assign empty_89_fu_567_p2 = zext_ln459_1_fu_557_p1 + 3'd1;
  assign grp_fu_309_p2 = word_q1 ^ statemt_q1;
  assign grp_fu_315_p2 = word_q0 ^ statemt_q0;
  assign grp_fu_321_p4 = { { statemt_q1[30:7] } };
  assign grp_fu_331_p4 = { { statemt_q0[30:7] } };
  assign icmp_ln447_fu_607_p2 = (and_ln_fu_599_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln451_fu_667_p2 = (and_ln1_fu_659_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln455_fu_725_p2 = (and_ln2_fu_717_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln460_fu_765_p2 = (and_ln3_fu_757_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln463_fu_803_p2 = (and_ln4_fu_795_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln467_fu_865_p2 = (and_ln5_fu_857_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln476_fu_933_p2 = (and_ln6_fu_925_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln480_fu_999_p2 = (and_ln7_fu_991_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln483_fu_1045_p2 = (and_ln8_fu_1037_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln489_fu_1085_p2 = (and_ln9_fu_1077_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln492_fu_1129_p2 = (and_ln10_fu_1121_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln495_fu_1175_p2 = (and_ln11_fu_1167_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln510_fu_371_p2 = (j_fu_82 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln519_fu_494_p2 = (j_4_fu_90 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln520_fu_531_p2 = (i_6_reg_298 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln531_fu_1227_p2 = (i_fu_94 == 3'd4)? 1'b1 : 1'b0;
  assign iv_rem_fu_573_p3 = (empty_88_fu_561_p2[0:0] == 1'b1)? 3'd0 : empty_89_fu_567_p2;
  assign mul_fu_351_p3 = { { n }, { 2'd0 } };
  assign or_ln1_fu_907_p3 = { { empty_86_reg_1373 }, { add_ln488_fu_902_p2 } };
  assign or_ln515_fu_425_p2 = shl_ln_fu_412_p3 | 4'd1;
  assign or_ln516_fu_471_p2 = ~(shl_ln_reg_1322 & ~4'd2);
  assign or_ln517_fu_481_p2 = shl_ln_reg_1322 | 4'd3;
  assign or_ln536_fu_1256_p2 = ~shl_ln1_fu_1243_p3 | 4'd1;
  assign or_ln537_fu_1272_p2 = ~shl_ln1_reg_1448 | 4'd2;
  assign or_ln538_fu_1282_p2 = ~shl_ln1_reg_1448 | 4'd3;
  assign or_ln_fu_890_p3 = { { empty_86_reg_1373 }, { xor_ln475_fu_885_p2 } };
  assign ret_d0 = xor_ln528_5_fu_1212_p2 ^ xor_ln528_2_fu_1200_p2;
  assign select_ln447_fu_631_p3 = (icmp_ln447_fu_607_p2[0:0] == 1'b1)? xor_ln447_fu_625_p2 : trunc_ln_fu_617_p3;
  assign select_ln451_fu_685_p3 = (icmp_ln451_fu_667_p2[0:0] == 1'b1)? xor_ln451_fu_679_p2 : shl_ln452_fu_673_p2;
  assign select_ln455_fu_737_p3 = (icmp_ln455_fu_725_p2[0:0] == 1'b1)? xor_ln456_fu_731_p2 : x_assign_2_fu_699_p3;
  assign select_ln460_fu_777_p3 = (icmp_ln460_fu_765_p2[0:0] == 1'b1)? xor_ln461_fu_771_p2 : trunc_ln1_fu_749_p3;
  assign select_ln463_fu_821_p3 = (icmp_ln463_fu_803_p2[0:0] == 1'b1)? xor_ln463_fu_815_p2 : shl_ln464_fu_809_p2;
  assign select_ln467_fu_877_p3 = (icmp_ln467_fu_865_p2[0:0] == 1'b1)? xor_ln468_fu_871_p2 : x_assign_8_fu_839_p3;
  assign select_ln476_fu_957_p3 = (icmp_ln476_fu_933_p2[0:0] == 1'b1)? xor_ln476_fu_951_p2 : trunc_ln2_fu_943_p3;
  assign select_ln480_fu_1011_p3 = (icmp_ln480_fu_999_p2[0:0] == 1'b1)? xor_ln481_fu_1005_p2 : shl_ln474_fu_975_p2;
  assign select_ln483_fu_1057_p3 = (icmp_ln483_fu_1045_p2[0:0] == 1'b1)? xor_ln484_fu_1051_p2 : x_assign_s_fu_1019_p3;
  assign select_ln489_fu_1097_p3 = (icmp_ln489_fu_1085_p2[0:0] == 1'b1)? xor_ln490_fu_1091_p2 : trunc_ln474_1_fu_1069_p3;
  assign select_ln492_fu_1141_p3 = (icmp_ln492_fu_1129_p2[0:0] == 1'b1)? xor_ln493_fu_1135_p2 : shl_ln474_1_fu_1105_p2;
  assign select_ln495_fu_1187_p3 = (icmp_ln495_fu_1175_p2[0:0] == 1'b1)? xor_ln496_fu_1181_p2 : x_assign_1_fu_1149_p3;
  assign shl_ln1_fu_1243_p3 = { ~{ trunc_ln535_fu_1239_p1 }, ~{ 2'd0 } };
  assign shl_ln452_fu_673_p2 = xor_ln450_fu_643_p2 << 31'd1;
  assign shl_ln464_fu_809_p2 = select_ln460_fu_777_p3 << 31'd1;
  assign shl_ln474_1_fu_1105_p2 = select_ln489_fu_1097_p3 << 31'd1;
  assign shl_ln474_fu_975_p2 = xor_ln479_fu_969_p2 << 31'd1;
  assign shl_ln_fu_412_p3 = ~{ { ~trunc_ln514_fu_408_p1 }, { ~2'd0 } };
  assign tmp_21_fu_649_p4 = { { xor_ln450_fu_643_p2[30:7] } };
  assign tmp_22_fu_707_p4 = { { xor_ln454_fu_693_p2[30:7] } };
  assign tmp_24_fu_785_p4 = { { select_ln460_fu_777_p3[30:7] } };
  assign tmp_25_fu_847_p4 = { { xor_ln466_fu_833_p2[30:7] } };
  assign tmp_27_fu_981_p4 = { { xor_ln479_fu_969_p2[30:7] } };
  assign tmp_28_fu_1027_p4 = { { select_ln480_fu_1011_p3[30:7] } };
  assign tmp_30_fu_1111_p4 = { { select_ln489_fu_1097_p3[30:7] } };
  assign tmp_31_fu_1157_p4 = { { select_ln492_fu_1141_p3[30:7] } };
  assign tmp_s_fu_510_p3 = { { empty_86_fu_506_p1 }, { 2'd0 } };
  assign trunc_ln1_fu_749_p3 = { { trunc_ln445_fu_745_p1 }, { 1'd0 } };
  assign trunc_ln2_fu_943_p3 = { { trunc_ln477_fu_939_p1 }, { 1'd0 } };
  assign trunc_ln445_fu_745_p1 = statemt_q0[29:0];
  assign trunc_ln448_fu_613_p1 = statemt_q1[29:0];
  assign trunc_ln449_fu_639_p1 = statemt_q1[30:0];
  assign trunc_ln459_fu_553_p1 = i_6_reg_298[1:0];
  assign trunc_ln465_fu_829_p1 = statemt_q0[30:0];
  assign trunc_ln474_1_fu_1069_p3 = { { trunc_ln474_fu_1065_p1 }, { 1'd0 } };
  assign trunc_ln474_fu_1065_p1 = statemt_q0[29:0];
  assign trunc_ln477_fu_939_p1 = statemt_q1[29:0];
  assign trunc_ln478_fu_965_p1 = statemt_q1[30:0];
  assign trunc_ln514_fu_408_p1 = j_fu_82[1:0];
  assign trunc_ln535_fu_1239_p1 = i_fu_94[1:0];
  assign trunc_ln_fu_617_p3 = { { trunc_ln448_fu_613_p1 }, { 1'd0 } };
  assign x_assign_1_fu_1149_p3 = { { select_ln492_fu_1141_p3 }, { 1'd0 } };
  assign x_assign_2_fu_699_p3 = { { xor_ln454_fu_693_p2 }, { 1'd0 } };
  assign x_assign_8_fu_839_p3 = { ~(~{ ~xor_ln466_fu_833_p2 }), ~(~{ ~1'd0 }) };
  assign x_assign_s_fu_1019_p3 = { { select_ln480_fu_1011_p3 }, { 1'd0 } };
  assign xor_ln447_fu_625_p2 = trunc_ln_fu_617_p3 ^ 31'd283;
  assign xor_ln450_fu_643_p2 = trunc_ln449_fu_639_p1 ^ select_ln447_fu_631_p3;
  assign xor_ln451_fu_679_p2 = shl_ln452_fu_673_p2 ^ 31'd283;
  assign xor_ln454_fu_693_p2 = trunc_ln449_fu_639_p1 ^ select_ln451_fu_685_p3;
  assign xor_ln456_fu_731_p2 = x_assign_2_fu_699_p3 ^ 32'd283;
  assign xor_ln461_fu_771_p2 = trunc_ln1_fu_749_p3 ^ 31'd283;
  assign xor_ln463_fu_815_p2 = shl_ln464_fu_809_p2 ^ 31'd283;
  assign xor_ln466_fu_833_p2 = ~(~trunc_ln465_fu_829_p1 ^ select_ln463_fu_821_p3);
  assign xor_ln468_fu_871_p2 = ~(~x_assign_8_fu_839_p3) ^ 32'd283;
  assign xor_ln475_fu_885_p2 = trunc_ln459_reg_1414 ^ 2'd2;
  assign xor_ln476_fu_951_p2 = trunc_ln2_fu_943_p3 ^ 31'd283;
  assign xor_ln479_fu_969_p2 = trunc_ln478_fu_965_p1 ^ select_ln476_fu_957_p3;
  assign xor_ln481_fu_1005_p2 = shl_ln474_fu_975_p2 ^ 31'd283;
  assign xor_ln484_fu_1051_p2 = x_assign_s_fu_1019_p3 ^ 32'd283;
  assign xor_ln490_fu_1091_p2 = trunc_ln474_1_fu_1069_p3 ^ 31'd283;
  assign xor_ln493_fu_1135_p2 = shl_ln474_1_fu_1105_p2 ^ 31'd283;
  assign xor_ln496_fu_1181_p2 = x_assign_1_fu_1149_p3 ^ 32'd283;
  assign xor_ln528_1_fu_1195_p2 = statemt_q0 ^ ~statemt_load_29_reg_1425;
  assign xor_ln528_2_fu_1200_p2 = xor_ln528_1_fu_1195_p2 ^ statemt_q1;
  assign xor_ln528_3_fu_919_p2 = select_ln467_fu_877_p3 ^ select_ln455_fu_737_p3;
  assign xor_ln528_4_fu_1206_p2 = select_ln495_fu_1187_p3 ^ select_ln483_fu_1057_p3;
  assign xor_ln528_5_fu_1212_p2 = xor_ln528_4_fu_1206_p2 ^ ~xor_ln528_3_reg_1440;
  assign zext_ln446_fu_548_p1 = add_ln446_fu_543_p2;
  assign zext_ln459_1_fu_557_p1 = trunc_ln459_fu_553_p1;
  assign zext_ln459_2_fu_581_p1 = iv_rem_fu_573_p3;
  assign zext_ln459_fu_590_p1 = add_ln459_1_fu_585_p2;
  assign zext_ln475_fu_897_p1 = or_ln_fu_890_p3;
  assign zext_ln488_fu_914_p1 = or_ln1_fu_907_p3;
  assign zext_ln510_fu_367_p1 = j_fu_82;
  assign zext_ln514_1_fu_420_p1 = ~shl_ln_fu_412_p3;
  assign zext_ln514_2_fu_446_p1 = add_ln514_reg_1307;
  assign zext_ln514_3_fu_393_p1 = add_ln514_fu_383_p2;
  assign zext_ln514_fu_388_p1 = add_ln514_fu_383_p2;
  assign zext_ln515_1_fu_403_p1 = add_ln515_fu_397_p2;
  assign zext_ln515_fu_431_p1 = or_ln515_fu_425_p2;
  assign zext_ln516_1_fu_455_p1 = add_ln516_fu_449_p2;
  assign zext_ln516_fu_476_p1 = or_ln516_fu_471_p2;
  assign zext_ln517_1_fu_466_p1 = add_ln517_fu_460_p2;
  assign zext_ln517_fu_486_p1 = or_ln517_fu_481_p2;
  assign zext_ln520_1_fu_527_p1 = i_6_reg_298;
  assign zext_ln520_fu_518_p1 = tmp_s_fu_510_p3;
  assign zext_ln535_fu_1251_p1 = ~shl_ln1_fu_1243_p3;
  assign zext_ln536_fu_1262_p1 = or_ln536_fu_1256_p2;
  assign zext_ln537_fu_1277_p1 = or_ln537_fu_1272_p2;
  assign zext_ln538_fu_1287_p1 = or_ln538_fu_1282_p2;

  always @(posedge ap_clk) begin
    mul_reg_1299[1:0] <= 2'b00;
    shl_ln_reg_1322[1:0] <= 2'b00;
    statemt_addr_reg_1328[1:0] <= ~2'b00;
    statemt_addr_reg_1328[4] <= ~1'b0;
    statemt_addr_12_reg_1333[1:0] <= 2'b01;
    statemt_addr_12_reg_1333[4] <= 1'b0;
    statemt_addr_13_reg_1355[1:0] <= ~2'b10;
    statemt_addr_13_reg_1355[4] <= ~1'b0;
    statemt_addr_14_reg_1360[1:0] <= 2'b11;
    statemt_addr_14_reg_1360[4] <= 1'b0;
    tmp_s_reg_1379[1:0] <= 2'b00;
    zext_ln520_reg_1384[1:0] <= 2'b00;
    zext_ln520_reg_1384[4] <= 1'b0;
    zext_ln446_reg_1404[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    shl_ln1_reg_1448[1:0] <= ~2'b00;
    zext_ln535_reg_1454[1:0] <= 2'b00;
    zext_ln535_reg_1454[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    zext_ln536_reg_1464[1:0] <= 2'b01;
    zext_ln536_reg_1464[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    zext_ln537_reg_1474[1:0] <= 2'b10;
    zext_ln537_reg_1474[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    zext_ln538_reg_1484[1:0] <= 2'b11;
    zext_ln538_reg_1484[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
  end


endmodule


