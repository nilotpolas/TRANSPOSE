`timescale 1 ns / 1 ps


module aes_main_decrypt_1
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt_address0,
  statemt_ce0,
  statemt_we0,
  statemt_d0,
  statemt_q0,
  key_address0,
  key_ce0,
  key_q0
);

  parameter ap_ST_fsm_state1 = 28'd1;
  parameter ap_ST_fsm_state2 = 28'd2;
  parameter ap_ST_fsm_state3 = 28'd4;
  parameter ap_ST_fsm_state4 = 28'd8;
  parameter ap_ST_fsm_state5 = 28'd16;
  parameter ap_ST_fsm_state6 = 28'd32;
  parameter ap_ST_fsm_state7 = 28'd64;
  parameter ap_ST_fsm_state8 = 28'd128;
  parameter ap_ST_fsm_state9 = 28'd256;
  parameter ap_ST_fsm_state10 = 28'd512;
  parameter ap_ST_fsm_state11 = 28'd1024;
  parameter ap_ST_fsm_state12 = 28'd2048;
  parameter ap_ST_fsm_state13 = 28'd4096;
  parameter ap_ST_fsm_state14 = 28'd8192;
  parameter ap_ST_fsm_state15 = 28'd16384;
  parameter ap_ST_fsm_state16 = 28'd32768;
  parameter ap_ST_fsm_state17 = 28'd65536;
  parameter ap_ST_fsm_state18 = 28'd131072;
  parameter ap_ST_fsm_state19 = 28'd262144;
  parameter ap_ST_fsm_state20 = 28'd524288;
  parameter ap_ST_fsm_state21 = 28'd1048576;
  parameter ap_ST_fsm_state22 = 28'd2097152;
  parameter ap_ST_fsm_state23 = 28'd4194304;
  parameter ap_ST_fsm_state24 = 28'd8388608;
  parameter ap_ST_fsm_state25 = 28'd16777216;
  parameter ap_ST_fsm_state26 = 28'd33554432;
  parameter ap_ST_fsm_state27 = 28'd67108864;
  parameter ap_ST_fsm_state28 = 28'd134217728;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt_address0;
  output statemt_ce0;
  output statemt_we0;
  output [31:0] statemt_d0;
  input [31:0] statemt_q0;
  output [4:0] key_address0;
  output key_ce0;
  input [7:0] key_q0;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg key_ce0;
  (* fsm_encoding = "none" *)
  reg [27:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  reg [8:0] word_address0;
  reg word_ce0;
  reg word_we0;
  reg [31:0] word_d0;
  wire [31:0] word_q0;
  reg [8:0] word_address1;
  reg word_ce1;
  wire [31:0] word_q1;
  wire [7:0] Sbox_address0;
  reg Sbox_ce0;
  wire [7:0] Sbox_q0;
  wire [7:0] Sbox_address1;
  reg Sbox_ce1;
  wire [7:0] Sbox_q1;
  wire [7:0] Sbox_address2;
  reg Sbox_ce2;
  wire [7:0] Sbox_q2;
  wire [7:0] Sbox_address3;
  reg Sbox_ce3;
  wire [7:0] Sbox_q3;
  wire [4:0] Rcon0_address0;
  reg Rcon0_ce0;
  wire [7:0] Rcon0_q0;
  reg [4:0] statemt_r_address0;
  reg statemt_r_ce0;
  reg statemt_r_we0;
  reg [31:0] statemt_r_d0;
  wire [31:0] statemt_r_q0;
  reg [4:0] statemt_r_address1;
  reg statemt_r_ce1;
  reg statemt_r_we1;
  reg [31:0] statemt_r_d1;
  wire [31:0] statemt_r_q1;
  wire [31:0] grp_fu_577_p2;
  reg [31:0] reg_589;
  wire ap_CS_fsm_state16;
  wire ap_CS_fsm_state24;
  wire ap_CS_fsm_state25;
  wire [31:0] grp_fu_583_p2;
  reg [31:0] reg_594;
  wire [2:0] add_ln71_fu_613_p2;
  reg [2:0] add_ln71_reg_1782;
  wire ap_CS_fsm_state2;
  wire [3:0] tmp_2_fu_623_p3;
  reg [3:0] tmp_2_reg_1787;
  wire [0:0] icmp_ln71_fu_607_p2;
  reg [8:0] word_addr_4_reg_1799;
  wire ap_CS_fsm_state3;
  wire [2:0] add_ln75_fu_698_p2;
  reg [2:0] add_ln75_reg_1807;
  wire [0:0] icmp_ln75_fu_692_p2;
  wire [8:0] zext_ln83_fu_726_p1;
  reg [8:0] zext_ln83_reg_1820;
  wire ap_CS_fsm_state5;
  wire [5:0] add_ln90_fu_736_p2;
  reg [5:0] add_ln90_reg_1828;
  wire [0:0] icmp_ln83_fu_730_p2;
  wire [8:0] zext_ln90_3_fu_742_p1;
  reg [8:0] zext_ln90_3_reg_1833;
  wire ap_CS_fsm_state6;
  reg [31:0] temp_1_1_reg_1865;
  wire [3:0] trunc_ln98_fu_791_p1;
  reg [3:0] trunc_ln98_reg_1872;
  wire [7:0] trunc_ln98_1_fu_795_p1;
  reg [7:0] trunc_ln98_1_reg_1878;
  reg [31:0] temp_2_1_reg_1883;
  wire [3:0] trunc_ln99_fu_799_p1;
  reg [3:0] trunc_ln99_reg_1890;
  wire [7:0] trunc_ln99_1_fu_803_p1;
  reg [7:0] trunc_ln99_1_reg_1896;
  wire ap_CS_fsm_state7;
  wire [0:0] icmp_ln88_fu_810_p2;
  wire [31:0] zext_ln90_2_fu_1308_p1;
  wire ap_CS_fsm_state8;
  wire [31:0] zext_ln91_fu_1312_p1;
  wire [31:0] zext_ln92_fu_1316_p1;
  wire [31:0] zext_ln95_fu_1320_p1;
  wire [8:0] zext_ln110_fu_1329_p1;
  reg [8:0] zext_ln110_reg_1959;
  wire ap_CS_fsm_state9;
  wire ap_CS_fsm_state10;
  reg [8:0] word_addr_10_reg_1969;
  wire [2:0] add_ln110_fu_1389_p2;
  reg [2:0] add_ln110_reg_1977;
  wire [31:0] tmp_fu_1395_p6;
  reg [31:0] tmp_reg_1982;
  wire [0:0] icmp_ln110_fu_1383_p2;
  wire [63:0] zext_ln11_fu_1428_p1;
  reg [63:0] zext_ln11_reg_1987;
  wire ap_CS_fsm_state12;
  wire [0:0] icmp_ln11_fu_1433_p2;
  wire [5:0] zext_ln570_cast_fu_1470_p3;
  reg [5:0] zext_ln570_cast_reg_2010;
  wire ap_CS_fsm_state14;
  wire [0:0] icmp_ln566_fu_1458_p2;
  wire [3:0] shl_ln_fu_1502_p3;
  reg [3:0] shl_ln_reg_2025;
  reg [4:0] statemt_addr_2_reg_2031;
  reg [4:0] statemt_addr_3_reg_2037;
  wire ap_CS_fsm_state15;
  wire [31:0] xor_ln570_fu_1561_p2;
  reg [31:0] xor_ln570_reg_2060;
  wire [31:0] xor_ln571_fu_1567_p2;
  reg [31:0] xor_ln571_reg_2065;
  reg [4:0] statemt_addr_4_reg_2070;
  reg [4:0] statemt_addr_5_reg_2075;
  reg [3:0] i_7_reg_2080;
  wire ap_CS_fsm_state19;
  wire ap_CS_fsm_state23;
  reg [8:0] word_addr_13_reg_2105;
  reg [8:0] word_addr_14_reg_2110;
  wire [3:0] shl_ln570_1_fu_1690_p3;
  reg [3:0] shl_ln570_1_reg_2118;
  wire [0:0] icmp_ln566_1_fu_1674_p2;
  reg [4:0] statemt_addr_6_reg_2124;
  reg [4:0] statemt_addr_7_reg_2129;
  reg [4:0] statemt_addr_8_reg_2141;
  reg [4:0] statemt_addr_9_reg_2146;
  wire [63:0] zext_ln34_fu_1747_p1;
  reg [63:0] zext_ln34_reg_2151;
  wire ap_CS_fsm_state27;
  wire [0:0] icmp_ln34_fu_1752_p2;
  wire grp_InversShiftRow_ByteSub_fu_560_ap_start;
  wire grp_InversShiftRow_ByteSub_fu_560_ap_done;
  wire grp_InversShiftRow_ByteSub_fu_560_ap_idle;
  wire grp_InversShiftRow_ByteSub_fu_560_ap_ready;
  wire [4:0] grp_InversShiftRow_ByteSub_fu_560_statemt_address0;
  wire grp_InversShiftRow_ByteSub_fu_560_statemt_ce0;
  wire grp_InversShiftRow_ByteSub_fu_560_statemt_we0;
  wire [31:0] grp_InversShiftRow_ByteSub_fu_560_statemt_d0;
  wire [4:0] grp_InversShiftRow_ByteSub_fu_560_statemt_address1;
  wire grp_InversShiftRow_ByteSub_fu_560_statemt_ce1;
  wire grp_InversShiftRow_ByteSub_fu_560_statemt_we1;
  wire [31:0] grp_InversShiftRow_ByteSub_fu_560_statemt_d1;
  wire grp_AddRoundKey_InversMixColumn_fu_568_ap_start;
  wire grp_AddRoundKey_InversMixColumn_fu_568_ap_done;
  wire grp_AddRoundKey_InversMixColumn_fu_568_ap_idle;
  wire grp_AddRoundKey_InversMixColumn_fu_568_ap_ready;
  wire [8:0] grp_AddRoundKey_InversMixColumn_fu_568_word_address0;
  wire grp_AddRoundKey_InversMixColumn_fu_568_word_ce0;
  wire [8:0] grp_AddRoundKey_InversMixColumn_fu_568_word_address1;
  wire grp_AddRoundKey_InversMixColumn_fu_568_word_ce1;
  wire [4:0] grp_AddRoundKey_InversMixColumn_fu_568_statemt_address0;
  wire grp_AddRoundKey_InversMixColumn_fu_568_statemt_ce0;
  wire grp_AddRoundKey_InversMixColumn_fu_568_statemt_we0;
  wire [31:0] grp_AddRoundKey_InversMixColumn_fu_568_statemt_d0;
  wire [4:0] grp_AddRoundKey_InversMixColumn_fu_568_statemt_address1;
  wire grp_AddRoundKey_InversMixColumn_fu_568_statemt_ce1;
  wire grp_AddRoundKey_InversMixColumn_fu_568_statemt_we1;
  wire [31:0] grp_AddRoundKey_InversMixColumn_fu_568_statemt_d1;
  reg [2:0] i_reg_498;
  wire ap_CS_fsm_state4;
  reg [31:0] temp_2_0_reg_509;
  reg [31:0] temp_1_0_reg_519;
  reg [31:0] temp_0_0_reg_529;
  reg [31:0] temp_3_reg_539;
  reg [2:0] i_2_reg_549;
  wire ap_CS_fsm_state11;
  reg grp_InversShiftRow_ByteSub_fu_560_ap_start_reg;
  wire ap_CS_fsm_state21;
  wire ap_CS_fsm_state18;
  wire ap_CS_fsm_state22;
  reg grp_AddRoundKey_InversMixColumn_fu_568_ap_start_reg;
  wire [0:0] icmp_ln25_fu_1597_p2;
  wire ap_CS_fsm_state20;
  wire [63:0] zext_ln79_4_fu_683_p1;
  wire [63:0] zext_ln79_fu_709_p1;
  wire [63:0] zext_ln90_5_fu_756_p1;
  wire [63:0] zext_ln91_1_fu_767_p1;
  wire [63:0] zext_ln92_1_fu_786_p1;
  wire [63:0] zext_ln90_1_fu_777_p1;
  wire [63:0] zext_ln216_2_fu_937_p1;
  wire [63:0] zext_ln90_fu_957_p1;
  wire [63:0] zext_ln216_5_fu_1067_p1;
  wire [63:0] zext_ln216_8_fu_1182_p1;
  wire [63:0] zext_ln216_11_fu_1297_p1;
  wire [63:0] zext_ln114_1_fu_1368_p1;
  wire [63:0] zext_ln114_2_fu_1378_p1;
  wire ap_CS_fsm_state13;
  wire [63:0] zext_ln570_fu_1478_p1;
  wire [63:0] zext_ln571_2_fu_1493_p1;
  wire [63:0] zext_ln570_1_fu_1510_p1;
  wire [63:0] zext_ln571_fu_1521_p1;
  wire [63:0] zext_ln572_2_fu_1545_p1;
  wire [63:0] zext_ln573_2_fu_1556_p1;
  wire [63:0] zext_ln572_fu_1578_p1;
  wire [63:0] zext_ln573_fu_1588_p1;
  wire [63:0] zext_ln566_fu_1622_p1;
  wire [63:0] zext_ln571_3_fu_1639_p1;
  wire [63:0] zext_ln572_3_fu_1656_p1;
  wire [63:0] zext_ln573_3_fu_1669_p1;
  wire [63:0] zext_ln570_2_fu_1698_p1;
  wire [63:0] zext_ln571_1_fu_1709_p1;
  wire [63:0] zext_ln572_1_fu_1729_p1;
  wire [63:0] zext_ln573_1_fu_1739_p1;
  wire ap_CS_fsm_state28;
  reg [2:0] j_fu_158;
  reg [5:0] j_1_fu_162;
  wire [5:0] add_ln83_fu_1409_p2;
  reg [5:0] i_1_fu_166;
  wire [5:0] add_ln11_fu_1439_p2;
  reg [2:0] j_2_fu_170;
  wire [2:0] add_ln566_fu_1464_p2;
  reg [3:0] i_3_fu_174;
  wire [3:0] i_8_fu_1603_p2;
  reg [2:0] j_3_fu_178;
  wire [2:0] add_ln566_1_fu_1680_p2;
  reg [5:0] i_5_fu_182;
  wire [5:0] add_ln34_fu_1758_p2;
  wire [31:0] zext_ln79_1_fu_718_p1;
  wire [31:0] xor_ln114_fu_1419_p2;
  wire ap_CS_fsm_state17;
  wire ap_CS_fsm_state26;
  wire [1:0] empty_27_fu_619_p1;
  wire [9:0] tmp_3_fu_636_p3;
  wire [5:0] tmp_4_fu_648_p3;
  wire [10:0] zext_ln79_2_fu_644_p1;
  wire [10:0] zext_ln79_3_fu_656_p1;
  wire [10:0] sub_ln79_fu_660_p2;
  wire [5:0] tmp_6_cast_fu_666_p4;
  wire [8:0] tmp_7_fu_676_p3;
  wire [3:0] zext_ln75_fu_688_p1;
  wire [3:0] add_ln79_fu_704_p2;
  wire [7:0] zext_ln90_4_fu_746_p1;
  wire [7:0] add_ln90_2_fu_750_p2;
  wire [8:0] add_ln91_fu_761_p2;
  wire [8:0] add_ln92_fu_781_p2;
  wire [1:0] empty_30_fu_807_p1;
  wire [7:0] sub_ln216_fu_839_p2;
  wire [3:0] trunc_ln216_4_fu_844_p4;
  wire [0:0] tmp_1_fu_832_p3;
  wire [3:0] sub_ln216_1_fu_854_p2;
  wire [3:0] tmp_8_fu_860_p4;
  wire [3:0] select_ln216_fu_869_p3;
  wire [4:0] p_and_f1_fu_885_p3;
  wire [3:0] sub_ln216_8_fu_896_p2;
  wire [4:0] p_and_t1_fu_901_p3;
  wire [5:0] zext_ln216_1_fu_909_p1;
  wire [5:0] sub_ln216_9_fu_913_p2;
  wire [5:0] zext_ln216_fu_892_p1;
  wire [5:0] select_ln216_1_fu_919_p3;
  wire [7:0] tmp_9_fu_877_p3;
  wire signed [7:0] sext_ln216_fu_927_p1;
  wire [7:0] add_ln216_fu_931_p2;
  wire [3:0] trunc_ln5_fu_942_p4;
  wire [3:0] add_ln90_1_fu_951_p2;
  wire [7:0] sub_ln216_2_fu_969_p2;
  wire [3:0] trunc_ln216_6_fu_974_p4;
  wire [0:0] tmp_5_fu_962_p3;
  wire [3:0] sub_ln216_3_fu_984_p2;
  wire [3:0] tmp_s_fu_990_p4;
  wire [3:0] select_ln216_2_fu_999_p3;
  wire [4:0] p_and_f2_fu_1015_p3;
  wire [3:0] sub_ln216_10_fu_1026_p2;
  wire [4:0] p_and_t2_fu_1031_p3;
  wire [5:0] zext_ln216_4_fu_1039_p1;
  wire [5:0] sub_ln216_11_fu_1043_p2;
  wire [5:0] zext_ln216_3_fu_1022_p1;
  wire [5:0] select_ln216_3_fu_1049_p3;
  wire [7:0] tmp_6_fu_1007_p3;
  wire signed [7:0] sext_ln216_1_fu_1057_p1;
  wire [7:0] add_ln216_1_fu_1061_p2;
  wire [7:0] trunc_ln93_1_fu_820_p1;
  wire [7:0] sub_ln216_4_fu_1080_p2;
  wire [3:0] trunc_ln216_8_fu_1086_p4;
  wire [0:0] tmp_10_fu_1072_p3;
  wire [3:0] sub_ln216_5_fu_1096_p2;
  wire [3:0] tmp_11_fu_1102_p4;
  wire [3:0] select_ln216_4_fu_1112_p3;
  wire [3:0] trunc_ln93_fu_816_p1;
  wire [4:0] p_and_f4_fu_1128_p3;
  wire [3:0] sub_ln216_12_fu_1140_p2;
  wire [4:0] p_and_t6_fu_1146_p3;
  wire [5:0] zext_ln216_7_fu_1154_p1;
  wire [5:0] sub_ln216_13_fu_1158_p2;
  wire [5:0] zext_ln216_6_fu_1136_p1;
  wire [5:0] select_ln216_5_fu_1164_p3;
  wire [7:0] tmp_12_fu_1120_p3;
  wire signed [7:0] sext_ln216_2_fu_1172_p1;
  wire [7:0] add_ln216_2_fu_1176_p2;
  wire [7:0] trunc_ln97_1_fu_828_p1;
  wire [7:0] sub_ln216_6_fu_1195_p2;
  wire [3:0] trunc_ln216_s_fu_1201_p4;
  wire [0:0] tmp_13_fu_1187_p3;
  wire [3:0] sub_ln216_7_fu_1211_p2;
  wire [3:0] tmp_14_fu_1217_p4;
  wire [3:0] select_ln216_6_fu_1227_p3;
  wire [3:0] trunc_ln97_fu_824_p1;
  wire [4:0] p_and_f_fu_1243_p3;
  wire [3:0] sub_ln216_14_fu_1255_p2;
  wire [4:0] p_and_t_fu_1261_p3;
  wire [5:0] zext_ln216_10_fu_1269_p1;
  wire [5:0] sub_ln216_15_fu_1273_p2;
  wire [5:0] zext_ln216_9_fu_1251_p1;
  wire [5:0] select_ln216_7_fu_1279_p3;
  wire [7:0] tmp_15_fu_1235_p3;
  wire signed [7:0] sext_ln216_3_fu_1287_p1;
  wire [7:0] add_ln216_3_fu_1291_p2;
  wire [7:0] temp_0_1_fu_1302_p2;
  wire [5:0] empty_31_fu_1324_p2;
  wire [1:0] trunc_ln114_fu_1333_p1;
  wire [5:0] tmp_17_fu_1345_p3;
  wire [8:0] tmp_16_fu_1337_p3;
  wire [8:0] zext_ln114_fu_1353_p1;
  wire [8:0] sub_ln114_fu_1357_p2;
  wire [8:0] add_ln114_fu_1363_p2;
  wire [8:0] add_ln114_1_fu_1373_p2;
  wire [7:0] zext_ln570_4_fu_1483_p1;
  wire [7:0] add_ln571_fu_1487_p2;
  wire [1:0] trunc_ln570_fu_1498_p1;
  wire [3:0] or_ln571_fu_1515_p2;
  wire [8:0] zext_ln570_3_fu_1536_p1;
  wire [8:0] add_ln572_fu_1539_p2;
  wire [8:0] add_ln573_fu_1550_p2;
  wire [3:0] or_ln572_fu_1573_p2;
  wire [3:0] or_ln573_fu_1583_p2;
  wire [3:0] tmp_18_fu_1627_p3;
  wire signed [6:0] sext_ln571_fu_1635_p1;
  wire [4:0] tmp_19_fu_1644_p3;
  wire signed [7:0] sext_ln572_fu_1652_p1;
  wire [8:0] tmp_29_cast_fu_1661_p3;
  wire [1:0] trunc_ln570_1_fu_1686_p1;
  wire [3:0] or_ln571_1_fu_1703_p2;
  wire [3:0] or_ln572_1_fu_1724_p2;
  wire [3:0] or_ln573_1_fu_1734_p2;
  reg [27:0] ap_NS_fsm;
  reg ap_ST_fsm_state1_blk;
  wire ap_ST_fsm_state2_blk;
  wire ap_ST_fsm_state3_blk;
  wire ap_ST_fsm_state4_blk;
  wire ap_ST_fsm_state5_blk;
  wire ap_ST_fsm_state6_blk;
  wire ap_ST_fsm_state7_blk;
  wire ap_ST_fsm_state8_blk;
  wire ap_ST_fsm_state9_blk;
  wire ap_ST_fsm_state10_blk;
  wire ap_ST_fsm_state11_blk;
  wire ap_ST_fsm_state12_blk;
  wire ap_ST_fsm_state13_blk;
  wire ap_ST_fsm_state14_blk;
  wire ap_ST_fsm_state15_blk;
  wire ap_ST_fsm_state16_blk;
  wire ap_ST_fsm_state17_blk;
  reg ap_ST_fsm_state18_blk;
  wire ap_ST_fsm_state19_blk;
  reg ap_ST_fsm_state20_blk;
  wire ap_ST_fsm_state21_blk;
  reg ap_ST_fsm_state22_blk;
  wire ap_ST_fsm_state23_blk;
  wire ap_ST_fsm_state24_blk;
  wire ap_ST_fsm_state25_blk;
  wire ap_ST_fsm_state26_blk;
  wire ap_ST_fsm_state27_blk;
  wire ap_ST_fsm_state28_blk;
  wire ap_ce_reg;

  initial begin
    #0 ap_CS_fsm = 28'd1;
    #0 grp_InversShiftRow_ByteSub_fu_560_ap_start_reg = 1'b0;
    #0 grp_AddRoundKey_InversMixColumn_fu_568_ap_start_reg = 1'b0;
  end


  aes_main_decrypt_1_word_RAM_AUTO_1R1W
  #(
    .DataWidth(32),
    .AddressRange(480),
    .AddressWidth(9)
  )
  word_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(word_address0),
    .ce0(word_ce0),
    .we0(word_we0),
    .d0(word_d0),
    .q0(word_q0),
    .address1(word_address1),
    .ce1(word_ce1),
    .q1(word_q1)
  );


  aes_main_decrypt_1_Sbox_ROM_AUTO_1R
  #(
    .DataWidth(8),
    .AddressRange(256),
    .AddressWidth(8)
  )
  Sbox_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(Sbox_address0),
    .ce0(Sbox_ce0),
    .q0(Sbox_q0),
    .address1(Sbox_address1),
    .ce1(Sbox_ce1),
    .q1(Sbox_q1),
    .address2(Sbox_address2),
    .ce2(Sbox_ce2),
    .q2(Sbox_q2),
    .address3(Sbox_address3),
    .ce3(Sbox_ce3),
    .q3(Sbox_q3)
  );


  aes_main_decrypt_1_Rcon0_ROM_AUTO_1R
  #(
    .DataWidth(8),
    .AddressRange(30),
    .AddressWidth(5)
  )
  Rcon0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(Rcon0_address0),
    .ce0(Rcon0_ce0),
    .q0(Rcon0_q0)
  );


  aes_main_decrypt_1_statemt_r_RAM_AUTO_1R1W
  #(
    .DataWidth(32),
    .AddressRange(32),
    .AddressWidth(5)
  )
  statemt_r_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(statemt_r_address0),
    .ce0(statemt_r_ce0),
    .we0(statemt_r_we0),
    .d0(statemt_r_d0),
    .q0(statemt_r_q0),
    .address1(statemt_r_address1),
    .ce1(statemt_r_ce1),
    .we1(statemt_r_we1),
    .d1(~statemt_r_d1),
    .q1(statemt_r_q1)
  );


  aes_main_InversShiftRow_ByteSub
  grp_InversShiftRow_ByteSub_fu_560
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_InversShiftRow_ByteSub_fu_560_ap_start),
    .ap_done(grp_InversShiftRow_ByteSub_fu_560_ap_done),
    .ap_idle(grp_InversShiftRow_ByteSub_fu_560_ap_idle),
    .ap_ready(grp_InversShiftRow_ByteSub_fu_560_ap_ready),
    .statemt_address0(grp_InversShiftRow_ByteSub_fu_560_statemt_address0),
    .statemt_ce0(grp_InversShiftRow_ByteSub_fu_560_statemt_ce0),
    .statemt_we0(grp_InversShiftRow_ByteSub_fu_560_statemt_we0),
    .statemt_d0(grp_InversShiftRow_ByteSub_fu_560_statemt_d0),
    .statemt_q0(statemt_r_q0),
    .statemt_address1(grp_InversShiftRow_ByteSub_fu_560_statemt_address1),
    .statemt_ce1(grp_InversShiftRow_ByteSub_fu_560_statemt_ce1),
    .statemt_we1(grp_InversShiftRow_ByteSub_fu_560_statemt_we1),
    .statemt_d1(grp_InversShiftRow_ByteSub_fu_560_statemt_d1),
    .statemt_q1(statemt_r_q1)
  );


  aes_main_AddRoundKey_InversMixColumn
  grp_AddRoundKey_InversMixColumn_fu_568
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_AddRoundKey_InversMixColumn_fu_568_ap_start),
    .ap_done(grp_AddRoundKey_InversMixColumn_fu_568_ap_done),
    .ap_idle(grp_AddRoundKey_InversMixColumn_fu_568_ap_idle),
    .ap_ready(grp_AddRoundKey_InversMixColumn_fu_568_ap_ready),
    .n(i_7_reg_2080),
    .word_address0(grp_AddRoundKey_InversMixColumn_fu_568_word_address0),
    .word_ce0(grp_AddRoundKey_InversMixColumn_fu_568_word_ce0),
    .word_q0(word_q0),
    .word_address1(grp_AddRoundKey_InversMixColumn_fu_568_word_address1),
    .word_ce1(grp_AddRoundKey_InversMixColumn_fu_568_word_ce1),
    .word_q1(word_q1),
    .statemt_address0(grp_AddRoundKey_InversMixColumn_fu_568_statemt_address0),
    .statemt_ce0(grp_AddRoundKey_InversMixColumn_fu_568_statemt_ce0),
    .statemt_we0(grp_AddRoundKey_InversMixColumn_fu_568_statemt_we0),
    .statemt_d0(grp_AddRoundKey_InversMixColumn_fu_568_statemt_d0),
    .statemt_q0(statemt_r_q0),
    .statemt_address1(grp_AddRoundKey_InversMixColumn_fu_568_statemt_address1),
    .statemt_ce1(grp_AddRoundKey_InversMixColumn_fu_568_statemt_ce1),
    .statemt_we1(grp_AddRoundKey_InversMixColumn_fu_568_statemt_we1),
    .statemt_d1(grp_AddRoundKey_InversMixColumn_fu_568_statemt_d1),
    .statemt_q1(statemt_r_q1)
  );


  aes_main_mux_42_32_1_1
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(32),
    .din1_WIDTH(32),
    .din2_WIDTH(32),
    .din3_WIDTH(32),
    .din4_WIDTH(2),
    .dout_WIDTH(32)
  )
  mux_42_32_1_1_U7
  (
    .din0(temp_0_0_reg_529),
    .din1(temp_1_0_reg_519),
    .din2(temp_2_0_reg_509),
    .din3(temp_3_reg_539),
    .din4(trunc_ln114_fu_1333_p1),
    .dout(tmp_fu_1395_p6)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_AddRoundKey_InversMixColumn_fu_568_ap_start_reg <= 1'b0;
    end else begin
      if((icmp_ln25_fu_1597_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state19)) begin
        grp_AddRoundKey_InversMixColumn_fu_568_ap_start_reg <= 1'b1;
      end else if(grp_AddRoundKey_InversMixColumn_fu_568_ap_ready == 1'b1) begin
        grp_AddRoundKey_InversMixColumn_fu_568_ap_start_reg <= 1'b0;
      end 
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_InversShiftRow_ByteSub_fu_560_ap_start_reg <= 1'b0;
    end else begin
      if((1'b1 == ap_CS_fsm_state21) | (icmp_ln566_fu_1458_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state14)) begin
        grp_InversShiftRow_ByteSub_fu_560_ap_start_reg <= 1'b1;
      end else if(grp_InversShiftRow_ByteSub_fu_560_ap_ready == 1'b1) begin
        grp_InversShiftRow_ByteSub_fu_560_ap_start_reg <= 1'b0;
      end 
    end
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state5) & (icmp_ln83_fu_730_p2 == 1'd1)) begin
      i_1_fu_166 <= 6'd0;
    end else if((icmp_ln11_fu_1433_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state12)) begin
      i_1_fu_166 <= add_ln11_fu_1439_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      i_2_reg_549 <= 3'd0;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      i_2_reg_549 <= add_ln110_reg_1977;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln566_fu_1458_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state14)) begin
      i_3_fu_174 <= 4'd9;
    end else if((icmp_ln25_fu_1597_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state19)) begin
      i_3_fu_174 <= i_8_fu_1603_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln566_1_fu_1674_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state23)) begin
      i_5_fu_182 <= 6'd0;
    end else if((icmp_ln34_fu_1752_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state27)) begin
      i_5_fu_182 <= add_ln34_fu_1758_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state2) & (icmp_ln71_fu_607_p2 == 1'd0)) begin
      i_reg_498 <= 3'd0;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      i_reg_498 <= add_ln75_reg_1807;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state2) & (icmp_ln71_fu_607_p2 == 1'd1)) begin
      j_1_fu_162 <= 6'd4;
    end else if((icmp_ln110_fu_1383_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state10)) begin
      j_1_fu_162 <= add_ln83_fu_1409_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln11_fu_1433_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state12)) begin
      j_2_fu_170 <= 3'd0;
    end else if((icmp_ln566_fu_1458_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      j_2_fu_170 <= add_ln566_fu_1464_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln25_fu_1597_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state19)) begin
      j_3_fu_178 <= 3'd0;
    end else if((icmp_ln566_1_fu_1674_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state23)) begin
      j_3_fu_178 <= add_ln566_1_fu_1680_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      j_fu_158 <= 3'd0;
    end else if((1'b1 == ap_CS_fsm_state3) & (icmp_ln75_fu_692_p2 == 1'd1)) begin
      j_fu_158 <= add_ln71_reg_1782;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln88_fu_810_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      temp_0_0_reg_529 <= word_q1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      temp_0_0_reg_529 <= zext_ln90_2_fu_1308_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln88_fu_810_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      temp_1_0_reg_519 <= ~temp_1_1_reg_1865;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      temp_1_0_reg_519 <= zext_ln91_fu_1312_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln88_fu_810_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      temp_2_0_reg_509 <= ~temp_2_1_reg_1883;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      temp_2_0_reg_509 <= zext_ln92_fu_1316_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln88_fu_810_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      temp_3_reg_539 <= word_q0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      temp_3_reg_539 <= zext_ln95_fu_1320_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      add_ln110_reg_1977 <= add_ln110_fu_1389_p2;
      word_addr_10_reg_1969 <= zext_ln114_2_fu_1378_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      add_ln71_reg_1782 <= add_ln71_fu_613_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      add_ln75_reg_1807 <= add_ln75_fu_698_p2;
      word_addr_4_reg_1799 <= zext_ln79_4_fu_683_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state5) & (icmp_ln83_fu_730_p2 == 1'd0)) begin
      add_ln90_reg_1828 <= add_ln90_fu_736_p2;
      zext_ln90_3_reg_1833[5:0] <= zext_ln90_3_fu_742_p1[5:0];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state19) begin
      i_7_reg_2080 <= i_3_fu_174;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state16)) begin
      reg_589 <= grp_fu_577_p2;
      reg_594 <= grp_fu_583_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln566_1_fu_1674_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state23)) begin
      shl_ln570_1_reg_2118[3:2] <= shl_ln570_1_fu_1690_p3[3:2];
      statemt_addr_6_reg_2124[3:2] <= zext_ln570_2_fu_1698_p1[3:2];
      statemt_addr_7_reg_2129[3:2] <= zext_ln571_1_fu_1709_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln566_fu_1458_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      shl_ln_reg_2025[3:2] <= shl_ln_fu_1502_p3[3:2];
      statemt_addr_2_reg_2031[3:2] <= zext_ln570_1_fu_1510_p1[3:2];
      statemt_addr_3_reg_2037[3:2] <= zext_ln571_fu_1521_p1[3:2];
      zext_ln570_cast_reg_2010[2:0] <= zext_ln570_cast_fu_1470_p3[2:0];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state15) begin
      statemt_addr_4_reg_2070[3:2] <= zext_ln572_fu_1578_p1[3:2];
      statemt_addr_5_reg_2075[3:2] <= zext_ln573_fu_1588_p1[3:2];
      xor_ln570_reg_2060 <= ~xor_ln570_fu_1561_p2;
      xor_ln571_reg_2065 <= ~xor_ln571_fu_1567_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state24) begin
      statemt_addr_8_reg_2141[3:2] <= zext_ln572_1_fu_1729_p1[3:2];
      statemt_addr_9_reg_2146[3:2] <= zext_ln573_1_fu_1739_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      temp_1_1_reg_1865 <= ~word_q1;
      temp_2_1_reg_1883 <= ~word_q0;
      trunc_ln98_1_reg_1878 <= trunc_ln98_1_fu_795_p1;
      trunc_ln98_reg_1872 <= trunc_ln98_fu_791_p1;
      trunc_ln99_1_reg_1896 <= trunc_ln99_1_fu_803_p1;
      trunc_ln99_reg_1890 <= trunc_ln99_fu_799_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state2) & (icmp_ln71_fu_607_p2 == 1'd0)) begin
      tmp_2_reg_1787[3:2] <= tmp_2_fu_623_p3[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln110_fu_1383_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state10)) begin
      tmp_reg_1982 <= tmp_fu_1395_p6;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      word_addr_13_reg_2105[2:0] <= zext_ln572_3_fu_1656_p1[2:0];
      word_addr_14_reg_2110[2:0] <= zext_ln573_3_fu_1669_p1[2:0];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      zext_ln110_reg_1959[5:0] <= zext_ln110_fu_1329_p1[5:0];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      zext_ln11_reg_1987[5:0] <= zext_ln11_fu_1428_p1[5:0];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      zext_ln34_reg_2151[5:0] <= zext_ln34_fu_1747_p1[5:0];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      zext_ln83_reg_1820[5:0] <= zext_ln83_fu_726_p1[5:0];
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      Rcon0_ce0 = 1'b1;
    end else begin
      Rcon0_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_ce0 = 1'b1;
    end else begin
      Sbox_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_ce1 = 1'b1;
    end else begin
      Sbox_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_ce2 = 1'b1;
    end else begin
      Sbox_ce2 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_ce3 = 1'b1;
    end else begin
      Sbox_ce3 = 1'b0;
    end
  end

  assign ap_ST_fsm_state10_blk = 1'b0;
  assign ap_ST_fsm_state11_blk = 1'b0;
  assign ap_ST_fsm_state12_blk = 1'b0;
  assign ap_ST_fsm_state13_blk = 1'b0;
  assign ap_ST_fsm_state14_blk = 1'b0;
  assign ap_ST_fsm_state15_blk = 1'b0;
  assign ap_ST_fsm_state16_blk = 1'b0;
  assign ap_ST_fsm_state17_blk = 1'b0;

  always @(*) begin
    if(grp_InversShiftRow_ByteSub_fu_560_ap_done == 1'b0) begin
      ap_ST_fsm_state18_blk = 1'b1;
    end else begin
      ap_ST_fsm_state18_blk = 1'b0;
    end
  end

  assign ap_ST_fsm_state19_blk = 1'b0;

  always @(*) begin
    if(ap_start == 1'b0) begin
      ap_ST_fsm_state1_blk = 1'b1;
    end else begin
      ap_ST_fsm_state1_blk = 1'b0;
    end
  end


  always @(*) begin
    if(grp_AddRoundKey_InversMixColumn_fu_568_ap_done == 1'b0) begin
      ap_ST_fsm_state20_blk = 1'b1;
    end else begin
      ap_ST_fsm_state20_blk = 1'b0;
    end
  end

  assign ap_ST_fsm_state21_blk = 1'b0;

  always @(*) begin
    if(grp_InversShiftRow_ByteSub_fu_560_ap_done == 1'b0) begin
      ap_ST_fsm_state22_blk = 1'b1;
    end else begin
      ap_ST_fsm_state22_blk = 1'b0;
    end
  end

  assign ap_ST_fsm_state23_blk = 1'b0;
  assign ap_ST_fsm_state24_blk = 1'b0;
  assign ap_ST_fsm_state25_blk = 1'b0;
  assign ap_ST_fsm_state26_blk = 1'b0;
  assign ap_ST_fsm_state27_blk = 1'b0;
  assign ap_ST_fsm_state28_blk = 1'b0;
  assign ap_ST_fsm_state2_blk = 1'b0;
  assign ap_ST_fsm_state3_blk = 1'b0;
  assign ap_ST_fsm_state4_blk = 1'b0;
  assign ap_ST_fsm_state5_blk = 1'b0;
  assign ap_ST_fsm_state6_blk = 1'b0;
  assign ap_ST_fsm_state7_blk = 1'b0;
  assign ap_ST_fsm_state8_blk = 1'b0;
  assign ap_ST_fsm_state9_blk = 1'b0;

  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1) | (icmp_ln34_fu_1752_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state27)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((icmp_ln34_fu_1752_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state27)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      key_ce0 = 1'b1;
    end else begin
      key_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state28) begin
      statemt_address0 = zext_ln34_reg_2151;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address0 = zext_ln11_fu_1428_p1;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state12)) begin
      statemt_ce0 = 1'b1;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state26) begin
      statemt_r_address0 = statemt_addr_8_reg_2141;
    end else if(1'b1 == ap_CS_fsm_state25) begin
      statemt_r_address0 = statemt_addr_6_reg_2124;
    end else if(1'b1 == ap_CS_fsm_state24) begin
      statemt_r_address0 = zext_ln572_1_fu_1729_p1;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      statemt_r_address0 = zext_ln570_2_fu_1698_p1;
    end else if(1'b1 == ap_CS_fsm_state17) begin
      statemt_r_address0 = statemt_addr_4_reg_2070;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt_r_address0 = statemt_addr_2_reg_2031;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_r_address0 = zext_ln572_fu_1578_p1;
    end else if((icmp_ln566_fu_1458_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      statemt_r_address0 = zext_ln571_fu_1521_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_r_address0 = zext_ln11_reg_1987;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_address0 = grp_AddRoundKey_InversMixColumn_fu_568_statemt_address0;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_address0 = grp_InversShiftRow_ByteSub_fu_560_statemt_address0;
    end else begin
      statemt_r_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      statemt_r_address1 = zext_ln34_fu_1747_p1;
    end else if(1'b1 == ap_CS_fsm_state26) begin
      statemt_r_address1 = statemt_addr_9_reg_2146;
    end else if(1'b1 == ap_CS_fsm_state25) begin
      statemt_r_address1 = statemt_addr_7_reg_2129;
    end else if(1'b1 == ap_CS_fsm_state24) begin
      statemt_r_address1 = zext_ln573_1_fu_1739_p1;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      statemt_r_address1 = zext_ln571_1_fu_1709_p1;
    end else if(1'b1 == ap_CS_fsm_state17) begin
      statemt_r_address1 = statemt_addr_5_reg_2075;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt_r_address1 = statemt_addr_3_reg_2037;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_r_address1 = zext_ln573_fu_1588_p1;
    end else if((icmp_ln566_fu_1458_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      statemt_r_address1 = zext_ln570_1_fu_1510_p1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_address1 = grp_AddRoundKey_InversMixColumn_fu_568_statemt_address1;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_address1 = grp_InversShiftRow_ByteSub_fu_560_statemt_address1;
    end else begin
      statemt_r_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state16) | (icmp_ln566_fu_1458_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      statemt_r_ce0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_ce0 = grp_AddRoundKey_InversMixColumn_fu_568_statemt_ce0;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_ce0 = grp_InversShiftRow_ByteSub_fu_560_statemt_ce0;
    end else begin
      statemt_r_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state16) | (icmp_ln566_fu_1458_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      statemt_r_ce1 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_ce1 = grp_AddRoundKey_InversMixColumn_fu_568_statemt_ce1;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_ce1 = grp_InversShiftRow_ByteSub_fu_560_statemt_ce1;
    end else begin
      statemt_r_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state25)) begin
      statemt_r_d0 = reg_589;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt_r_d0 = ~xor_ln570_reg_2060;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_r_d0 = statemt_q0;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_d0 = grp_AddRoundKey_InversMixColumn_fu_568_statemt_d0;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_d0 = grp_InversShiftRow_ByteSub_fu_560_statemt_d0;
    end else begin
      statemt_r_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state25)) begin
      statemt_r_d1 = ~reg_594;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt_r_d1 = xor_ln571_reg_2065;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_d1 = ~grp_AddRoundKey_InversMixColumn_fu_568_statemt_d1;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_d1 = ~grp_InversShiftRow_ByteSub_fu_560_statemt_d1;
    end else begin
      statemt_r_d1 = ~'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state16)) begin
      statemt_r_we0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_we0 = grp_AddRoundKey_InversMixColumn_fu_568_statemt_we0;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_we0 = grp_InversShiftRow_ByteSub_fu_560_statemt_we0;
    end else begin
      statemt_r_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state16)) begin
      statemt_r_we1 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_r_we1 = grp_AddRoundKey_InversMixColumn_fu_568_statemt_we1;
    end else if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state18)) begin
      statemt_r_we1 = grp_InversShiftRow_ByteSub_fu_560_statemt_we1;
    end else begin
      statemt_r_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state28) begin
      statemt_we0 = 1'b1;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state24) begin
      word_address0 = word_addr_13_reg_2105;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      word_address0 = zext_ln566_fu_1622_p1;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      word_address0 = zext_ln572_2_fu_1545_p1;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      word_address0 = zext_ln570_fu_1478_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      word_address0 = word_addr_10_reg_1969;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      word_address0 = zext_ln92_1_fu_786_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      word_address0 = zext_ln91_1_fu_767_p1;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      word_address0 = word_addr_4_reg_1799;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      word_address0 = grp_AddRoundKey_InversMixColumn_fu_568_word_address0;
    end else begin
      word_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state24) begin
      word_address1 = word_addr_14_reg_2110;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      word_address1 = zext_ln571_3_fu_1639_p1;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      word_address1 = zext_ln573_2_fu_1556_p1;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      word_address1 = zext_ln571_2_fu_1493_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      word_address1 = zext_ln114_1_fu_1368_p1;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      word_address1 = zext_ln90_1_fu_777_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      word_address1 = zext_ln90_5_fu_756_p1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      word_address1 = grp_AddRoundKey_InversMixColumn_fu_568_word_address1;
    end else begin
      word_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state24)) begin
      word_ce0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      word_ce0 = grp_AddRoundKey_InversMixColumn_fu_568_word_ce0;
    end else begin
      word_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state24)) begin
      word_ce1 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      word_ce1 = grp_AddRoundKey_InversMixColumn_fu_568_word_ce1;
    end else begin
      word_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      word_d0 = xor_ln114_fu_1419_p2;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      word_d0 = zext_ln79_1_fu_718_p1;
    end else begin
      word_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      word_we0 = 1'b1;
    end else begin
      word_we0 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((1'b1 == ap_CS_fsm_state2) & (icmp_ln71_fu_607_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        if((1'b1 == ap_CS_fsm_state3) & (icmp_ln75_fu_692_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state3;
      end
      ap_ST_fsm_state5: begin
        if((1'b1 == ap_CS_fsm_state5) & (icmp_ln83_fu_730_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state6: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state7: begin
        if((icmp_ln88_fu_810_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        if((icmp_ln110_fu_1383_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state10)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state12: begin
        if((icmp_ln11_fu_1433_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state12)) begin
          ap_NS_fsm = ap_ST_fsm_state14;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state14: begin
        if((icmp_ln566_fu_1458_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state14)) begin
          ap_NS_fsm = ap_ST_fsm_state18;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state15;
        end
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state17: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state18: begin
        if((grp_InversShiftRow_ByteSub_fu_560_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state18)) begin
          ap_NS_fsm = ap_ST_fsm_state19;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state18;
        end
      end
      ap_ST_fsm_state19: begin
        if((icmp_ln25_fu_1597_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state19)) begin
          ap_NS_fsm = ap_ST_fsm_state23;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state20;
        end
      end
      ap_ST_fsm_state20: begin
        if((grp_AddRoundKey_InversMixColumn_fu_568_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state20)) begin
          ap_NS_fsm = ap_ST_fsm_state21;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state20;
        end
      end
      ap_ST_fsm_state21: begin
        ap_NS_fsm = ap_ST_fsm_state22;
      end
      ap_ST_fsm_state22: begin
        if((grp_InversShiftRow_ByteSub_fu_560_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state22)) begin
          ap_NS_fsm = ap_ST_fsm_state19;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state22;
        end
      end
      ap_ST_fsm_state23: begin
        if((icmp_ln566_1_fu_1674_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state23)) begin
          ap_NS_fsm = ap_ST_fsm_state27;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state24;
        end
      end
      ap_ST_fsm_state24: begin
        ap_NS_fsm = ap_ST_fsm_state25;
      end
      ap_ST_fsm_state25: begin
        ap_NS_fsm = ap_ST_fsm_state26;
      end
      ap_ST_fsm_state26: begin
        ap_NS_fsm = ap_ST_fsm_state23;
      end
      ap_ST_fsm_state27: begin
        if((icmp_ln34_fu_1752_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state27)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state28;
        end
      end
      ap_ST_fsm_state28: begin
        ap_NS_fsm = ap_ST_fsm_state27;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign Rcon0_address0 = zext_ln90_fu_957_p1;
  assign Sbox_address0 = zext_ln216_11_fu_1297_p1;
  assign Sbox_address1 = zext_ln216_8_fu_1182_p1;
  assign Sbox_address2 = zext_ln216_5_fu_1067_p1;
  assign Sbox_address3 = zext_ln216_2_fu_937_p1;
  assign add_ln110_fu_1389_p2 = i_2_reg_549 + 3'd1;
  assign add_ln114_1_fu_1373_p2 = sub_ln114_fu_1357_p2 + zext_ln83_reg_1820;
  assign add_ln114_fu_1363_p2 = sub_ln114_fu_1357_p2 + zext_ln110_reg_1959;
  assign add_ln11_fu_1439_p2 = i_1_fu_166 + 6'd1;
  assign add_ln216_1_fu_1061_p2 = $signed(tmp_6_fu_1007_p3) + $signed(sext_ln216_1_fu_1057_p1);
  assign add_ln216_2_fu_1176_p2 = $signed(tmp_12_fu_1120_p3) + $signed(sext_ln216_2_fu_1172_p1);
  assign add_ln216_3_fu_1291_p2 = $signed(tmp_15_fu_1235_p3) + $signed(sext_ln216_3_fu_1287_p1);
  assign add_ln216_fu_931_p2 = $signed(tmp_9_fu_877_p3) + $signed(sext_ln216_fu_927_p1);
  assign add_ln34_fu_1758_p2 = i_5_fu_182 + 6'd1;
  assign add_ln566_1_fu_1680_p2 = j_3_fu_178 + 3'd1;
  assign add_ln566_fu_1464_p2 = j_2_fu_170 + 3'd1;
  assign add_ln571_fu_1487_p2 = zext_ln570_4_fu_1483_p1 + 8'd120;
  assign add_ln572_fu_1539_p2 = zext_ln570_3_fu_1536_p1 + 9'd240;
  assign add_ln573_fu_1550_p2 = $signed(zext_ln570_3_fu_1536_p1) + $signed(9'd360);
  assign add_ln71_fu_613_p2 = j_fu_158 + 3'd1;
  assign add_ln75_fu_698_p2 = i_reg_498 + 3'd1;
  assign add_ln79_fu_704_p2 = zext_ln75_fu_688_p1 + tmp_2_reg_1787;
  assign add_ln83_fu_1409_p2 = j_1_fu_162 + 6'd1;
  assign add_ln90_1_fu_951_p2 = $signed(trunc_ln5_fu_942_p4) + $signed(4'd15);
  assign add_ln90_2_fu_750_p2 = zext_ln90_4_fu_746_p1 + 8'd120;
  assign add_ln90_fu_736_p2 = $signed(j_1_fu_162) + $signed(6'd63);
  assign add_ln91_fu_761_p2 = zext_ln90_3_fu_742_p1 + 9'd240;
  assign add_ln92_fu_781_p2 = $signed(zext_ln90_3_reg_1833) + $signed(9'd360);
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];
  assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];
  assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];
  assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];
  assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];
  assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign empty_27_fu_619_p1 = j_fu_158[1:0];
  assign empty_30_fu_807_p1 = j_1_fu_162[1:0];
  assign empty_31_fu_1324_p2 = $signed(j_1_fu_162) + $signed(6'd60);
  assign grp_AddRoundKey_InversMixColumn_fu_568_ap_start = grp_AddRoundKey_InversMixColumn_fu_568_ap_start_reg;
  assign grp_InversShiftRow_ByteSub_fu_560_ap_start = grp_InversShiftRow_ByteSub_fu_560_ap_start_reg;
  assign grp_fu_577_p2 = word_q0 ^ statemt_r_q0;
  assign grp_fu_583_p2 = word_q1 ^ statemt_r_q1;
  assign i_8_fu_1603_p2 = $signed(i_3_fu_174) + $signed(4'd15);
  assign icmp_ln110_fu_1383_p2 = (i_2_reg_549 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln11_fu_1433_p2 = (i_1_fu_166 == 6'd32)? 1'b1 : 1'b0;
  assign icmp_ln25_fu_1597_p2 = (i_3_fu_174 == 4'd0)? 1'b1 : 1'b0;
  assign icmp_ln34_fu_1752_p2 = (i_5_fu_182 == 6'd32)? 1'b1 : 1'b0;
  assign icmp_ln566_1_fu_1674_p2 = (j_3_fu_178 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln566_fu_1458_p2 = (j_2_fu_170 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln71_fu_607_p2 = (j_fu_158 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln75_fu_692_p2 = (i_reg_498 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln83_fu_730_p2 = (j_1_fu_162 == 6'd44)? 1'b1 : 1'b0;
  assign icmp_ln88_fu_810_p2 = (empty_30_fu_807_p1 == 2'd0)? 1'b1 : 1'b0;
  assign key_address0 = zext_ln79_fu_709_p1;
  assign or_ln571_1_fu_1703_p2 = shl_ln570_1_fu_1690_p3 | 4'd1;
  assign or_ln571_fu_1515_p2 = shl_ln_fu_1502_p3 | 4'd1;
  assign or_ln572_1_fu_1724_p2 = shl_ln570_1_reg_2118 | 4'd2;
  assign or_ln572_fu_1573_p2 = shl_ln_reg_2025 | 4'd2;
  assign or_ln573_1_fu_1734_p2 = shl_ln570_1_reg_2118 | 4'd3;
  assign or_ln573_fu_1583_p2 = shl_ln_reg_2025 | 4'd3;
  assign p_and_f1_fu_885_p3 = { { 1'd0 }, { trunc_ln98_reg_1872 } };
  assign p_and_f2_fu_1015_p3 = { { 1'd0 }, { trunc_ln99_reg_1890 } };
  assign p_and_f4_fu_1128_p3 = { { 1'd0 }, { trunc_ln93_fu_816_p1 } };
  assign p_and_f_fu_1243_p3 = { { 1'd0 }, { trunc_ln97_fu_824_p1 } };
  assign p_and_t1_fu_901_p3 = { { 1'd0 }, { sub_ln216_8_fu_896_p2 } };
  assign p_and_t2_fu_1031_p3 = { { 1'd0 }, { sub_ln216_10_fu_1026_p2 } };
  assign p_and_t6_fu_1146_p3 = { { 1'd0 }, { sub_ln216_12_fu_1140_p2 } };
  assign p_and_t_fu_1261_p3 = { { 1'd0 }, { sub_ln216_14_fu_1255_p2 } };
  assign select_ln216_1_fu_919_p3 = (tmp_1_fu_832_p3[0:0] == 1'b1)? sub_ln216_9_fu_913_p2 : zext_ln216_fu_892_p1;
  assign select_ln216_2_fu_999_p3 = (tmp_5_fu_962_p3[0:0] == 1'b1)? sub_ln216_3_fu_984_p2 : tmp_s_fu_990_p4;
  assign select_ln216_3_fu_1049_p3 = (tmp_5_fu_962_p3[0:0] == 1'b1)? sub_ln216_11_fu_1043_p2 : zext_ln216_3_fu_1022_p1;
  assign select_ln216_4_fu_1112_p3 = (tmp_10_fu_1072_p3[0:0] == 1'b1)? sub_ln216_5_fu_1096_p2 : tmp_11_fu_1102_p4;
  assign select_ln216_5_fu_1164_p3 = (tmp_10_fu_1072_p3[0:0] == 1'b1)? sub_ln216_13_fu_1158_p2 : zext_ln216_6_fu_1136_p1;
  assign select_ln216_6_fu_1227_p3 = (tmp_13_fu_1187_p3[0:0] == 1'b1)? sub_ln216_7_fu_1211_p2 : tmp_14_fu_1217_p4;
  assign select_ln216_7_fu_1279_p3 = (tmp_13_fu_1187_p3[0:0] == 1'b1)? sub_ln216_15_fu_1273_p2 : zext_ln216_9_fu_1251_p1;
  assign select_ln216_fu_869_p3 = (tmp_1_fu_832_p3[0:0] == 1'b1)? sub_ln216_1_fu_854_p2 : tmp_8_fu_860_p4;
  assign sext_ln216_1_fu_1057_p1 = $signed(select_ln216_3_fu_1049_p3);
  assign sext_ln216_2_fu_1172_p1 = $signed(select_ln216_5_fu_1164_p3);
  assign sext_ln216_3_fu_1287_p1 = $signed(select_ln216_7_fu_1279_p3);
  assign sext_ln216_fu_927_p1 = $signed(select_ln216_1_fu_919_p3);
  assign sext_ln571_fu_1635_p1 = $signed(tmp_18_fu_1627_p3);
  assign sext_ln572_fu_1652_p1 = $signed(tmp_19_fu_1644_p3);
  assign shl_ln570_1_fu_1690_p3 = { { trunc_ln570_1_fu_1686_p1 }, { 2'd0 } };
  assign shl_ln_fu_1502_p3 = { { trunc_ln570_fu_1498_p1 }, { 2'd0 } };
  assign statemt_d0 = statemt_r_q1;
  assign sub_ln114_fu_1357_p2 = tmp_16_fu_1337_p3 - zext_ln114_fu_1353_p1;
  assign sub_ln216_10_fu_1026_p2 = 4'd0 - trunc_ln99_reg_1890;
  assign sub_ln216_11_fu_1043_p2 = 6'd0 - zext_ln216_4_fu_1039_p1;
  assign sub_ln216_12_fu_1140_p2 = 4'd0 - trunc_ln93_fu_816_p1;
  assign sub_ln216_13_fu_1158_p2 = 6'd0 - zext_ln216_7_fu_1154_p1;
  assign sub_ln216_14_fu_1255_p2 = 4'd0 - trunc_ln97_fu_824_p1;
  assign sub_ln216_15_fu_1273_p2 = 6'd0 - zext_ln216_10_fu_1269_p1;
  assign sub_ln216_1_fu_854_p2 = 4'd0 - trunc_ln216_4_fu_844_p4;
  assign sub_ln216_2_fu_969_p2 = 8'd0 - trunc_ln99_1_reg_1896;
  assign sub_ln216_3_fu_984_p2 = 4'd0 - trunc_ln216_6_fu_974_p4;
  assign sub_ln216_4_fu_1080_p2 = 8'd0 - trunc_ln93_1_fu_820_p1;
  assign sub_ln216_5_fu_1096_p2 = 4'd0 - trunc_ln216_8_fu_1086_p4;
  assign sub_ln216_6_fu_1195_p2 = 8'd0 - trunc_ln97_1_fu_828_p1;
  assign sub_ln216_7_fu_1211_p2 = 4'd0 - trunc_ln216_s_fu_1201_p4;
  assign sub_ln216_8_fu_896_p2 = 4'd0 - trunc_ln98_reg_1872;
  assign sub_ln216_9_fu_913_p2 = 6'd0 - zext_ln216_1_fu_909_p1;
  assign sub_ln216_fu_839_p2 = 8'd0 - trunc_ln98_1_reg_1878;
  assign sub_ln79_fu_660_p2 = zext_ln79_2_fu_644_p1 - zext_ln79_3_fu_656_p1;
  assign temp_0_1_fu_1302_p2 = Sbox_q3 ^ Rcon0_q0;
  assign tmp_10_fu_1072_p3 = word_q0[32'd31];
  assign tmp_11_fu_1102_p4 = { { word_q0[7:4] } };
  assign tmp_12_fu_1120_p3 = { { select_ln216_4_fu_1112_p3 }, { 4'd0 } };
  assign tmp_13_fu_1187_p3 = word_q1[32'd31];
  assign tmp_14_fu_1217_p4 = { { word_q1[7:4] } };
  assign tmp_15_fu_1235_p3 = { { select_ln216_6_fu_1227_p3 }, { 4'd0 } };
  assign tmp_16_fu_1337_p3 = { { trunc_ln114_fu_1333_p1 }, { 7'd0 } };
  assign tmp_17_fu_1345_p3 = { { i_2_reg_549 }, { 3'd0 } };
  assign tmp_18_fu_1627_p3 = { { 1'd1 }, { j_3_fu_178 } };
  assign tmp_19_fu_1644_p3 = { { 2'd2 }, { j_3_fu_178 } };
  assign tmp_1_fu_832_p3 = ~temp_1_1_reg_1865[32'd31];
  assign tmp_29_cast_fu_1661_p3 = { { 6'd45 }, { j_3_fu_178 } };
  assign tmp_2_fu_623_p3 = { { empty_27_fu_619_p1 }, { 2'd0 } };
  assign tmp_3_fu_636_p3 = { { i_reg_498 }, { 7'd0 } };
  assign tmp_4_fu_648_p3 = { { i_reg_498 }, { 3'd0 } };
  assign tmp_5_fu_962_p3 = ~temp_2_1_reg_1883[32'd31];
  assign tmp_6_cast_fu_666_p4 = { { sub_ln79_fu_660_p2[8:3] } };
  assign tmp_6_fu_1007_p3 = { { select_ln216_2_fu_999_p3 }, { 4'd0 } };
  assign tmp_7_fu_676_p3 = { { tmp_6_cast_fu_666_p4 }, { j_fu_158 } };
  assign tmp_8_fu_860_p4 = { { ~temp_1_1_reg_1865[7:4] } };
  assign tmp_9_fu_877_p3 = { { select_ln216_fu_869_p3 }, { 4'd0 } };
  assign tmp_s_fu_990_p4 = { { ~temp_2_1_reg_1883[7:4] } };
  assign trunc_ln114_fu_1333_p1 = i_2_reg_549[1:0];
  assign trunc_ln216_4_fu_844_p4 = { { sub_ln216_fu_839_p2[7:4] } };
  assign trunc_ln216_6_fu_974_p4 = { { sub_ln216_2_fu_969_p2[7:4] } };
  assign trunc_ln216_8_fu_1086_p4 = { { sub_ln216_4_fu_1080_p2[7:4] } };
  assign trunc_ln216_s_fu_1201_p4 = { { sub_ln216_6_fu_1195_p2[7:4] } };
  assign trunc_ln570_1_fu_1686_p1 = j_3_fu_178[1:0];
  assign trunc_ln570_fu_1498_p1 = j_2_fu_170[1:0];
  assign trunc_ln5_fu_942_p4 = { { j_1_fu_162[5:2] } };
  assign trunc_ln93_1_fu_820_p1 = word_q0[7:0];
  assign trunc_ln93_fu_816_p1 = word_q0[3:0];
  assign trunc_ln97_1_fu_828_p1 = word_q1[7:0];
  assign trunc_ln97_fu_824_p1 = word_q1[3:0];
  assign trunc_ln98_1_fu_795_p1 = word_q1[7:0];
  assign trunc_ln98_fu_791_p1 = word_q1[3:0];
  assign trunc_ln99_1_fu_803_p1 = word_q0[7:0];
  assign trunc_ln99_fu_799_p1 = word_q0[3:0];
  assign xor_ln114_fu_1419_p2 = word_q1 ^ tmp_reg_1982;
  assign xor_ln570_fu_1561_p2 = word_q0 ^ statemt_r_q1;
  assign xor_ln571_fu_1567_p2 = word_q1 ^ statemt_r_q0;
  assign zext_ln110_fu_1329_p1 = empty_31_fu_1324_p2;
  assign zext_ln114_1_fu_1368_p1 = add_ln114_fu_1363_p2;
  assign zext_ln114_2_fu_1378_p1 = add_ln114_1_fu_1373_p2;
  assign zext_ln114_fu_1353_p1 = tmp_17_fu_1345_p3;
  assign zext_ln11_fu_1428_p1 = i_1_fu_166;
  assign zext_ln216_10_fu_1269_p1 = p_and_t_fu_1261_p3;
  assign zext_ln216_11_fu_1297_p1 = add_ln216_3_fu_1291_p2;
  assign zext_ln216_1_fu_909_p1 = p_and_t1_fu_901_p3;
  assign zext_ln216_2_fu_937_p1 = add_ln216_fu_931_p2;
  assign zext_ln216_3_fu_1022_p1 = p_and_f2_fu_1015_p3;
  assign zext_ln216_4_fu_1039_p1 = p_and_t2_fu_1031_p3;
  assign zext_ln216_5_fu_1067_p1 = add_ln216_1_fu_1061_p2;
  assign zext_ln216_6_fu_1136_p1 = p_and_f4_fu_1128_p3;
  assign zext_ln216_7_fu_1154_p1 = p_and_t6_fu_1146_p3;
  assign zext_ln216_8_fu_1182_p1 = add_ln216_2_fu_1176_p2;
  assign zext_ln216_9_fu_1251_p1 = p_and_f_fu_1243_p3;
  assign zext_ln216_fu_892_p1 = p_and_f1_fu_885_p3;
  assign zext_ln34_fu_1747_p1 = i_5_fu_182;
  assign zext_ln566_fu_1622_p1 = j_3_fu_178;
  assign zext_ln570_1_fu_1510_p1 = shl_ln_fu_1502_p3;
  assign zext_ln570_2_fu_1698_p1 = shl_ln570_1_fu_1690_p3;
  assign zext_ln570_3_fu_1536_p1 = zext_ln570_cast_reg_2010;
  assign zext_ln570_4_fu_1483_p1 = zext_ln570_cast_fu_1470_p3;
  assign zext_ln570_cast_fu_1470_p3 = { { 3'd5 }, { j_2_fu_170 } };
  assign zext_ln570_fu_1478_p1 = zext_ln570_cast_fu_1470_p3;
  assign zext_ln571_1_fu_1709_p1 = or_ln571_1_fu_1703_p2;
  assign zext_ln571_2_fu_1493_p1 = add_ln571_fu_1487_p2;
  assign zext_ln571_3_fu_1639_p1 = $unsigned(sext_ln571_fu_1635_p1);
  assign zext_ln571_fu_1521_p1 = or_ln571_fu_1515_p2;
  assign zext_ln572_1_fu_1729_p1 = or_ln572_1_fu_1724_p2;
  assign zext_ln572_2_fu_1545_p1 = add_ln572_fu_1539_p2;
  assign zext_ln572_3_fu_1656_p1 = $unsigned(sext_ln572_fu_1652_p1);
  assign zext_ln572_fu_1578_p1 = or_ln572_fu_1573_p2;
  assign zext_ln573_1_fu_1739_p1 = or_ln573_1_fu_1734_p2;
  assign zext_ln573_2_fu_1556_p1 = add_ln573_fu_1550_p2;
  assign zext_ln573_3_fu_1669_p1 = tmp_29_cast_fu_1661_p3;
  assign zext_ln573_fu_1588_p1 = or_ln573_fu_1583_p2;
  assign zext_ln75_fu_688_p1 = i_reg_498;
  assign zext_ln79_1_fu_718_p1 = key_q0;
  assign zext_ln79_2_fu_644_p1 = tmp_3_fu_636_p3;
  assign zext_ln79_3_fu_656_p1 = tmp_4_fu_648_p3;
  assign zext_ln79_4_fu_683_p1 = tmp_7_fu_676_p3;
  assign zext_ln79_fu_709_p1 = add_ln79_fu_704_p2;
  assign zext_ln83_fu_726_p1 = j_1_fu_162;
  assign zext_ln90_1_fu_777_p1 = add_ln90_reg_1828;
  assign zext_ln90_2_fu_1308_p1 = temp_0_1_fu_1302_p2;
  assign zext_ln90_3_fu_742_p1 = add_ln90_fu_736_p2;
  assign zext_ln90_4_fu_746_p1 = add_ln90_fu_736_p2;
  assign zext_ln90_5_fu_756_p1 = add_ln90_2_fu_750_p2;
  assign zext_ln90_fu_957_p1 = add_ln90_1_fu_951_p2;
  assign zext_ln91_1_fu_767_p1 = add_ln91_fu_761_p2;
  assign zext_ln91_fu_1312_p1 = Sbox_q2;
  assign zext_ln92_1_fu_786_p1 = add_ln92_fu_781_p2;
  assign zext_ln92_fu_1316_p1 = Sbox_q1;
  assign zext_ln95_fu_1320_p1 = Sbox_q0;

  always @(posedge ap_clk) begin
    tmp_2_reg_1787[1:0] <= 2'b00;
    zext_ln83_reg_1820[8:6] <= 3'b000;
    zext_ln90_3_reg_1833[8:6] <= 3'b000;
    zext_ln110_reg_1959[8:6] <= 3'b000;
    zext_ln11_reg_1987[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
    zext_ln570_cast_reg_2010[5:3] <= 3'b101;
    shl_ln_reg_2025[1:0] <= 2'b00;
    statemt_addr_2_reg_2031[1:0] <= 2'b00;
    statemt_addr_2_reg_2031[4] <= 1'b0;
    statemt_addr_3_reg_2037[1:0] <= 2'b01;
    statemt_addr_3_reg_2037[4] <= 1'b0;
    statemt_addr_4_reg_2070[1:0] <= 2'b10;
    statemt_addr_4_reg_2070[4] <= 1'b0;
    statemt_addr_5_reg_2075[1:0] <= 2'b11;
    statemt_addr_5_reg_2075[4] <= 1'b0;
    word_addr_13_reg_2105[8:3] <= 6'b011110;
    word_addr_14_reg_2110[8:3] <= 6'b101101;
    shl_ln570_1_reg_2118[1:0] <= 2'b00;
    statemt_addr_6_reg_2124[1:0] <= 2'b00;
    statemt_addr_6_reg_2124[4] <= 1'b0;
    statemt_addr_7_reg_2129[1:0] <= 2'b01;
    statemt_addr_7_reg_2129[4] <= 1'b0;
    statemt_addr_8_reg_2141[1:0] <= 2'b10;
    statemt_addr_8_reg_2141[4] <= 1'b0;
    statemt_addr_9_reg_2146[1:0] <= 2'b11;
    statemt_addr_9_reg_2146[4] <= 1'b0;
    zext_ln34_reg_2151[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
  end


endmodule


