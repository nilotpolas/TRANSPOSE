

module sbox
(
  clk,
  t,
  dec_0,
  dec_1,
  dec_255,
  dec_169,
  dec_129,
  dec_9,
  dec_72,
  dec_242,
  dec_243,
  dec_152,
  dec_240,
  dec_4,
  dec_15,
  dec_12,
  dec_2,
  dec_3,
  dec_36,
  dec_220,
  dec_11,
  dec_158,
  dec_45,
  dec_88,
  dec_99,
  r,
  y
);

  reg [7:0] y_reg121;
  reg [7:0] y_reg122;
  reg [7:0] y_reg123;
  reg [7:0] y_reg124;
  reg [7:0] y_reg125;
  reg [7:0] y_reg126;
  reg [7:0] y_reg127;
  reg [7:0] y_reg128;
  reg [7:0] y_reg129;
  reg [7:0] y_reg130;
  reg [7:0] y_reg131;
  reg [7:0] y_reg132;
  reg [7:0] y_reg133;
  reg [7:0] y_reg134;
  reg [7:0] y_reg135;
  reg [7:0] y_reg136;
  reg [7:0] y_reg137;
  reg [7:0] y_reg138;
  reg [7:0] y_reg139;
  reg [7:0] y_reg140;
  reg [7:0] y_reg141;
  reg [7:0] y_reg142;
  reg [7:0] y_reg143;
  reg [7:0] y_reg144;
  reg [7:0] y_reg145;
  reg [7:0] y_reg146;
  reg [7:0] y_reg147;
  reg [7:0] y_reg148;
  reg [7:0] y_reg149;
  reg [7:0] y_reg150;
  reg [7:0] y_reg151;
  reg [7:0] y_reg152;
  reg [7:0] y_reg153;
  reg [7:0] y_reg154;
  reg [7:0] y_reg155;
  reg [7:0] y_reg156;
  reg [7:0] y_reg157;
  reg [7:0] y_reg158;
  reg [7:0] y_reg159;
  reg [7:0] y_reg160;
  reg [7:0] y_reg161;
  reg [7:0] y_reg162;
  reg [7:0] y_reg163;
  reg [7:0] y_reg164;
  reg [7:0] y_reg165;
  reg [7:0] y_reg166;
  reg [7:0] y_reg167;
  reg [7:0] y_reg168;
  reg [7:0] y_reg169;
  reg [7:0] y_reg170;
  reg [7:0] y_reg171;
  reg [7:0] y_reg172;
  reg [7:0] y_reg173;
  reg [7:0] y_reg174;
  reg [7:0] y_reg175;
  reg [7:0] y_reg176;
  reg [7:0] y_reg177;
  reg [7:0] y_reg178;
  reg [7:0] y_reg179;
  reg [7:0] y_reg180;
  reg [7:0] y_reg181;
  reg [7:0] y_reg182;
  reg [7:0] y_reg183;
  reg [7:0] y_reg184;
  reg [7:0] y_reg185;
  reg [7:0] y_reg186;
  reg [7:0] y_reg187;
  reg [7:0] y_reg188;
  reg [7:0] y_reg189;
  reg [7:0] y_reg190;
  reg [7:0] y_reg191;
  reg [7:0] y_reg192;
  reg [7:0] y_reg193;
  reg [7:0] y_reg194;
  reg [7:0] y_reg195;
  reg [7:0] y_reg196;
  reg [7:0] y_reg197;
  reg [7:0] y_reg198;
  reg [7:0] y_reg199;
  reg [7:0] y_reg200;
  reg [7:0] y_reg201;
  reg [7:0] y_reg202;
  reg [7:0] y_reg203;
  reg [7:0] y_reg204;
  reg [7:0] y_reg205;
  reg [7:0] y_reg206;
  reg [7:0] y_reg207;
  reg [7:0] y_reg208;
  reg [7:0] y_reg209;
  reg [7:0] y_reg210;
  reg [7:0] y_reg211;
  reg [7:0] y_reg212;
  reg [7:0] y_reg213;
  reg [7:0] y_reg214;
  reg [7:0] y_reg215;
  reg [7:0] y_reg216;
  reg [7:0] y_reg217;
  reg [7:0] y_reg218;
  reg [7:0] y_reg219;
  reg [7:0] y_reg220;
  reg [7:0] y_reg221;
  reg [7:0] y_reg222;
  reg [7:0] y_reg223;
  reg [7:0] y_reg224;
  reg [7:0] y_reg225;
  reg [7:0] y_reg226;
  reg [7:0] y_reg227;
  reg [7:0] y_reg228;
  reg [7:0] y_reg229;
  reg [7:0] y_reg230;
  reg [7:0] y_reg231;
  reg [7:0] y_reg232;
  reg [7:0] y_reg233;
  reg [7:0] y_reg234;
  reg [7:0] y_reg235;
  reg [7:0] y_reg236;
  reg [7:0] y_reg237;
  reg [7:0] y_reg238;
  reg [7:0] y_reg239;
  reg [7:0] y_reg240;
  reg [7:0] y_reg241;
  reg [7:0] y_reg242;
  reg [7:0] y_reg243;
  reg [7:0] y_reg244;
  reg [7:0] y_reg245;
  reg [7:0] y_reg246;
  reg [7:0] y_reg247;
  reg [7:0] y_reg248;
  reg [7:0] y_reg249;
  reg [7:0] y_reg250;
  reg [7:0] y_reg251;
  reg [7:0] y_reg252;
  reg [7:0] y_reg253;
  reg [7:0] y_reg254;
  reg [7:0] y_reg255;
  reg [7:0] y_reg256;
  reg [7:0] y_reg257;
  reg [7:0] y_reg258;
  reg [7:0] y_reg259;
  reg [7:0] y_reg260;
  reg [7:0] y_reg261;
  reg [7:0] y_reg262;
  reg [7:0] y_reg263;
  reg [7:0] y_reg264;
  reg [7:0] y_reg265;
  reg [7:0] y_reg266;
  reg [7:0] y_reg267;
  reg [7:0] y_reg268;
  reg [7:0] y_reg269;
  reg [7:0] y_reg270;
  reg [7:0] y_reg271;
  reg [7:0] y_reg272;
  reg [7:0] y_reg273;
  reg [7:0] y_reg274;
  reg [7:0] y_reg275;
  reg [7:0] y_reg276;
  reg [7:0] y_reg277;
  reg [7:0] y_reg278;
  reg [7:0] y_reg279;
  reg [7:0] y_reg280;
  reg [7:0] y_reg281;
  reg [7:0] y_reg282;
  reg [7:0] y_reg283;
  reg [7:0] y_reg284;
  reg [7:0] y_reg285;
  reg [7:0] y_reg286;
  reg [7:0] y_reg287;
  reg [7:0] y_reg288;
  reg [7:0] y_reg289;
  reg [7:0] y_reg290;
  reg [7:0] y_reg291;
  reg [7:0] y_reg292;
  reg [7:0] y_reg293;
  reg [7:0] y_reg294;
  reg [7:0] y_reg295;
  reg [7:0] y_reg296;
  reg [7:0] y_reg297;
  reg [7:0] y_reg298;
  reg [7:0] y_reg299;
  reg [7:0] y_reg300;
  reg [7:0] y_reg301;
  reg [7:0] y_reg302;
  reg [7:0] y_reg303;
  reg [7:0] y_reg304;
  reg [7:0] y_reg305;
  reg [7:0] y_reg306;
  reg [7:0] y_reg307;
  reg [7:0] y_reg308;
  reg [7:0] y_reg309;
  reg [7:0] y_reg310;
  reg [7:0] y_reg311;
  reg [7:0] y_reg312;
  reg [7:0] y_reg313;
  reg [7:0] y_reg314;
  reg [7:0] y_reg315;
  reg [7:0] y_reg316;
  reg [7:0] y_reg317;
  reg [7:0] y_reg318;
  reg [7:0] y_reg319;
  reg [7:0] y_reg320;
  reg [7:0] y_reg321;
  reg [7:0] y_reg322;
  reg [7:0] y_reg323;
  reg [7:0] y_reg324;
  reg [7:0] y_reg325;
  reg [7:0] y_reg326;
  reg [7:0] y_reg327;
  reg [7:0] y_reg328;
  reg [7:0] y_reg329;
  reg [7:0] y_reg330;
  reg [7:0] y_reg331;
  reg [7:0] y_reg332;
  reg [7:0] y_reg333;
  reg [7:0] y_reg334;
  reg [7:0] y_reg335;
  reg [7:0] y_reg336;
  reg [7:0] y_reg337;
  reg [7:0] y_reg338;
  reg [7:0] y_reg339;
  reg [7:0] y_reg340;
  reg [7:0] y_reg341;
  reg [7:0] y_reg342;
  reg [7:0] y_reg343;
  reg [7:0] y_reg344;
  reg [7:0] y_reg345;
  reg [7:0] y_reg346;
  reg [7:0] y_reg347;
  reg [7:0] y_reg348;
  reg [7:0] y_reg349;
  reg [7:0] y_reg350;
  reg [7:0] y_reg351;
  reg [7:0] y_reg352;
  reg [7:0] y_reg353;
  reg [7:0] y_reg354;
  reg [7:0] y_reg355;
  reg [7:0] y_reg356;
  reg [7:0] y_reg357;
  reg [7:0] y_reg358;
  reg [7:0] y_reg359;
  reg [7:0] y_reg360;
  reg [7:0] y_reg361;
  reg [7:0] y_reg362;
  reg [7:0] y_reg363;
  reg [7:0] y_reg364;
  reg [7:0] y_reg365;
  reg [7:0] y_reg366;
  reg [7:0] y_reg367;
  reg [7:0] y_reg368;
  reg [7:0] y_reg369;
  reg [7:0] y_reg370;
  reg [7:0] y_reg371;
  reg [7:0] y_reg372;
  reg [7:0] y_reg373;
  reg [7:0] y_reg374;
  reg [7:0] y_reg375;
  reg [7:0] y_reg376;
  reg [7:0] y_reg377;
  reg [7:0] y_reg378;
  reg [7:0] y_reg379;
  reg [7:0] y_reg380;
  reg [7:0] y_reg381;
  reg [7:0] y_reg382;
  reg [7:0] y_reg383;
  reg [7:0] y_reg384;
  reg [7:0] y_reg385;
  reg [7:0] y_reg386;
  reg [7:0] y_reg387;
  reg [7:0] y_reg388;
  reg [7:0] y_reg389;
  reg [7:0] y_reg390;
  reg [7:0] y_reg391;
  reg [7:0] y_reg392;
  reg [7:0] y_reg393;
  reg [7:0] y_reg394;
  reg [7:0] y_reg395;
  reg [7:0] y_reg396;
  reg [7:0] y_reg397;
  reg [7:0] y_reg398;
  reg [7:0] y_reg399;
  reg [7:0] y_reg400;
  reg [7:0] y_reg401;
  reg [7:0] y_reg402;
  reg [7:0] y_reg403;
  reg [7:0] y_reg404;
  reg [7:0] y_reg405;
  reg [7:0] y_reg406;
  reg [7:0] y_reg407;
  reg [7:0] y_reg408;
  reg [7:0] y_reg409;
  reg [7:0] y_reg410;
  reg [7:0] y_reg411;
  reg [7:0] y_reg412;
  reg [7:0] y_reg413;
  reg [7:0] y_reg414;
  reg [7:0] y_reg415;
  reg [7:0] y_reg416;
  reg [7:0] y_reg417;
  reg [7:0] y_reg418;
  reg [7:0] y_reg419;
  reg [7:0] y_reg420;
  reg [7:0] y_reg421;
  reg [7:0] y_reg422;
  reg [7:0] y_reg423;
  reg [7:0] y_reg424;
  reg [7:0] y_reg425;
  reg [7:0] y_reg426;
  reg [7:0] y_reg427;
  reg [7:0] y_reg428;
  reg [7:0] y_reg429;
  reg [7:0] y_reg430;
  reg [7:0] y_reg431;
  reg [7:0] y_reg432;
  reg [7:0] y_reg433;
  reg [7:0] y_reg434;
  reg [7:0] y_reg435;
  reg [7:0] y_reg436;
  reg [7:0] y_reg437;
  reg [7:0] y_reg438;
  reg [7:0] y_reg439;
  reg [7:0] y_reg440;
  reg [7:0] y_reg441;
  reg [7:0] y_reg442;
  reg [7:0] y_reg443;
  reg [7:0] y_reg444;
  reg [7:0] y_reg445;
  reg [7:0] y_reg446;
  reg [7:0] y_reg447;
  reg [7:0] y_reg448;
  reg [7:0] y_reg449;
  reg [7:0] y_reg450;
  reg [7:0] y_reg451;
  reg [7:0] y_reg452;
  reg [7:0] y_reg453;
  reg [7:0] y_reg454;
  reg [7:0] y_reg455;
  reg [7:0] y_reg456;
  reg [7:0] y_reg457;
  reg [7:0] y_reg458;
  reg [7:0] y_reg459;
  reg [7:0] y_reg460;
  reg [7:0] y_reg461;
  reg [7:0] y_reg462;
  reg [7:0] y_reg463;
  reg [7:0] y_reg464;
  reg [7:0] y_reg465;
  reg [7:0] y_reg466;
  reg [7:0] y_reg467;
  reg [7:0] y_reg468;
  reg [7:0] y_reg469;
  reg [7:0] y_reg470;
  reg [7:0] y_reg471;
  reg [7:0] y_reg472;
  reg [7:0] y_reg473;
  reg [7:0] y_reg474;
  reg [7:0] y_reg475;
  reg [7:0] y_reg476;
  reg [7:0] y_reg477;
  reg [7:0] y_reg478;
  reg [7:0] y_reg479;
  reg [7:0] y_reg480;
  reg [7:0] y_reg481;
  reg [7:0] y_reg482;
  reg [7:0] y_reg483;
  reg [7:0] y_reg484;
  reg [7:0] y_reg485;
  reg [7:0] y_reg486;
  reg [7:0] y_reg487;
  reg [7:0] y_reg488;
  reg [7:0] y_reg489;
  reg [7:0] y_reg490;
  reg [7:0] y_reg491;
  reg [7:0] y_reg492;
  reg [7:0] y_reg493;
  reg [7:0] y_reg494;
  reg [7:0] y_reg495;
  reg [7:0] y_reg496;
  reg [7:0] y_reg497;
  reg [7:0] y_reg498;
  reg [7:0] y_reg499;
  reg [7:0] y_reg500;
  reg [7:0] y_reg501;
  reg [7:0] y_reg502;
  reg [7:0] y_reg503;
  reg [7:0] y_reg504;
  reg [7:0] y_reg505;
  reg [7:0] y_reg506;
  reg [7:0] y_reg507;
  reg [7:0] y_reg508;
  reg [7:0] y_reg509;
  reg [7:0] y_reg510;
  reg [7:0] y_reg511;
  reg [7:0] y_reg512;
  reg [7:0] y_reg513;
  reg [7:0] y_reg514;
  reg [7:0] y_reg515;
  reg [7:0] y_reg516;
  reg [7:0] y_reg517;
  reg [7:0] y_reg518;
  reg [7:0] y_reg519;
  reg [7:0] y_reg520;
  reg [7:0] y_reg521;
  reg [7:0] y_reg522;
  reg [7:0] y_reg523;
  reg [7:0] y_reg524;
  reg [7:0] y_reg525;
  reg [7:0] y_reg526;
  reg [7:0] y_reg527;
  reg [7:0] y_reg528;
  reg [7:0] y_reg529;
  reg [7:0] y_reg530;
  reg [7:0] y_reg531;
  reg [7:0] y_reg532;
  reg [7:0] y_reg533;
  reg [7:0] y_reg534;
  reg [7:0] y_reg535;
  reg [7:0] y_reg536;
  reg [7:0] y_reg537;
  reg [7:0] y_reg538;
  reg [7:0] y_reg539;
  reg [7:0] y_reg540;
  reg [7:0] y_reg541;
  reg [7:0] y_reg542;
  reg [7:0] y_reg543;
  reg [7:0] y_reg544;
  reg [7:0] y_reg545;
  reg [7:0] y_reg546;
  reg [7:0] y_reg547;
  reg [7:0] y_reg548;
  reg [7:0] y_reg549;
  reg [7:0] y_reg550;
  reg [7:0] y_reg551;
  reg [7:0] y_reg552;
  reg [7:0] y_reg553;
  reg [7:0] y_reg554;
  reg [7:0] y_reg555;
  reg [7:0] y_reg556;
  reg [7:0] y_reg557;
  reg [7:0] y_reg558;
  reg [7:0] y_reg559;
  reg [7:0] y_reg560;
  reg [7:0] y_reg561;
  reg [7:0] y_reg562;
  reg [7:0] y_reg563;
  reg [7:0] y_reg564;
  reg [7:0] y_reg565;
  reg [7:0] y_reg566;
  reg [7:0] y_reg567;
  reg [7:0] y_reg568;
  reg [7:0] y_reg569;
  reg [7:0] y_reg570;
  reg [7:0] y_reg571;
  reg [7:0] y_reg572;
  reg [7:0] y_reg573;
  reg [7:0] y_reg574;
  reg [7:0] y_reg575;
  reg [7:0] y_reg576;
  reg [7:0] y_reg577;
  reg [7:0] y_reg578;
  reg [7:0] y_reg579;
  reg [7:0] y_reg580;
  reg [7:0] y_reg581;
  reg [7:0] y_reg582;
  reg [7:0] y_reg583;
  reg [7:0] y_reg584;
  reg [7:0] y_reg585;
  reg [7:0] y_reg586;
  reg [7:0] y_reg587;
  reg [7:0] y_reg588;
  reg [7:0] y_reg589;
  reg [7:0] y_reg590;
  reg [7:0] y_reg591;
  reg [7:0] y_reg592;
  reg [7:0] y_reg593;
  reg [7:0] y_reg594;
  reg [7:0] y_reg595;
  reg [7:0] y_reg596;
  reg [7:0] y_reg597;
  reg [7:0] y_reg598;
  reg [7:0] y_reg599;
  reg [7:0] y_reg600;
  reg [7:0] y_reg601;
  reg [7:0] y_reg602;
  reg [7:0] y_reg603;
  reg [7:0] y_reg604;
  reg [7:0] y_reg605;
  reg [7:0] y_reg606;
  reg [7:0] y_reg607;
  reg [7:0] y_reg608;
  reg [7:0] y_reg609;
  reg [7:0] y_reg610;
  reg [7:0] y_reg611;
  reg [7:0] y_reg612;
  reg [7:0] y_reg613;
  reg [7:0] y_reg614;
  reg [7:0] y_reg615;
  reg [7:0] y_reg616;
  reg [7:0] y_reg617;
  reg [7:0] y_reg618;
  reg [7:0] y_reg619;
  reg [7:0] y_reg620;
  reg [7:0] y_reg621;
  reg [7:0] y_reg622;
  reg [7:0] y_reg623;
  reg [7:0] y_reg624;
  reg [7:0] y_reg625;
  reg [7:0] y_reg626;
  reg [7:0] y_reg627;
  reg [7:0] y_reg628;
  reg [7:0] y_reg629;
  reg [7:0] y_reg630;
  reg [7:0] y_reg631;
  reg [7:0] y_reg632;
  reg [7:0] y_reg633;
  reg [7:0] y_reg634;
  reg [7:0] y_reg635;
  reg [7:0] y_reg636;
  reg [7:0] y_reg637;
  reg [7:0] y_reg638;
  reg [7:0] y_reg639;
  reg [7:0] y_reg640;
  reg [7:0] y_reg641;
  reg [7:0] y_reg642;
  reg [7:0] y_reg643;
  reg [7:0] y_reg644;
  reg [7:0] y_reg645;
  reg [7:0] y_reg646;
  reg [7:0] y_reg647;
  reg [7:0] y_reg648;
  reg [7:0] y_reg649;
  reg [7:0] y_reg650;
  reg [7:0] y_reg651;
  reg [7:0] y_reg652;
  reg [7:0] y_reg653;
  reg [7:0] y_reg654;
  reg [7:0] y_reg655;
  reg [7:0] y_reg656;
  reg [7:0] y_reg657;
  reg [7:0] y_reg658;
  reg [7:0] y_reg659;
  reg [7:0] y_reg660;
  reg [7:0] y_reg661;
  reg [7:0] y_reg662;
  reg [7:0] y_reg663;
  reg [7:0] y_reg664;
  reg [7:0] y_reg665;
  reg [7:0] y_reg666;
  reg [7:0] y_reg667;
  reg [7:0] y_reg668;
  reg [7:0] y_reg669;
  reg [7:0] y_reg670;
  reg [7:0] y_reg671;
  reg [7:0] y_reg672;
  reg [7:0] y_reg673;
  reg [7:0] y_reg674;
  reg [7:0] y_reg675;
  reg [7:0] y_reg676;
  reg [7:0] y_reg677;
  reg [7:0] y_reg678;
  reg [7:0] y_reg679;
  reg [7:0] y_reg680;
  reg [7:0] y_reg681;
  reg [7:0] y_reg682;
  reg [7:0] y_reg683;
  reg [7:0] y_reg684;
  reg [7:0] y_reg685;
  reg [7:0] y_reg686;
  reg [7:0] y_reg687;
  reg [7:0] y_reg688;
  reg [7:0] y_reg689;
  reg [7:0] y_reg690;
  reg [7:0] y_reg691;
  reg [7:0] y_reg692;
  reg [7:0] y_reg693;
  reg [7:0] y_reg694;
  reg [7:0] y_reg695;
  reg [7:0] y_reg696;
  reg [7:0] y_reg697;
  reg [7:0] y_reg698;
  reg [7:0] y_reg699;
  reg [7:0] y_reg700;
  reg [7:0] y_reg701;
  reg [7:0] y_reg702;
  reg [7:0] y_reg703;
  reg [7:0] y_reg704;
  reg [7:0] y_reg705;
  reg [7:0] y_reg706;
  reg [7:0] y_reg707;
  reg [7:0] y_reg708;
  reg [7:0] y_reg709;
  reg [7:0] y_reg710;
  reg [7:0] y_reg711;
  reg [7:0] y_reg712;
  reg [7:0] y_reg713;
  reg [7:0] y_reg714;
  reg [7:0] y_reg715;
  reg [7:0] y_reg716;
  reg [7:0] y_reg717;
  reg [7:0] y_reg718;
  reg [7:0] y_reg719;
  reg [7:0] y_reg720;
  reg [7:0] y_reg721;
  reg [7:0] y_reg722;
  reg [7:0] y_reg723;
  reg [7:0] y_reg724;
  reg [7:0] y_reg725;
  reg [7:0] y_reg726;
  reg [7:0] y_reg727;
  reg [7:0] y_reg728;
  reg [7:0] y_reg729;
  reg [7:0] y_reg730;
  reg [7:0] y_reg731;
  reg [7:0] y_reg732;
  reg [7:0] y_reg733;
  reg [7:0] y_reg734;
  reg [7:0] y_reg735;
  reg [7:0] y_reg736;
  reg [7:0] y_reg737;
  reg [7:0] y_reg738;
  reg [7:0] y_reg739;
  reg [7:0] y_reg740;
  reg [7:0] y_reg741;
  reg [7:0] y_reg742;
  reg [7:0] y_reg743;
  reg [7:0] y_reg744;
  reg [7:0] y_reg745;
  reg [7:0] y_reg746;
  reg [7:0] y_reg747;
  reg [7:0] y_reg748;
  reg [7:0] y_reg749;
  reg [7:0] y_reg750;
  reg [7:0] y_reg751;
  reg [7:0] y_reg752;
  reg [7:0] y_reg753;
  reg [7:0] y_reg754;
  reg [7:0] y_reg755;
  reg [7:0] y_reg756;
  reg [7:0] y_reg757;
  reg [7:0] y_reg758;
  reg [7:0] y_reg759;
  reg [7:0] y_reg760;
  reg [7:0] y_reg761;
  reg [7:0] y_reg762;
  reg [7:0] y_reg763;
  reg [7:0] y_reg764;
  reg [7:0] y_reg765;
  reg [7:0] y_reg766;
  reg [7:0] y_reg767;
  reg [7:0] y_reg768;
  reg [7:0] y_reg769;
  reg [7:0] y_reg770;
  reg [7:0] y_reg771;
  reg [7:0] y_reg772;
  reg [7:0] y_reg773;
  reg [7:0] y_reg774;
  reg [7:0] y_reg775;
  reg [7:0] y_reg776;
  reg [7:0] y_reg777;
  reg [7:0] y_reg778;
  reg [7:0] y_reg779;
  reg [7:0] y_reg780;
  reg [7:0] y_reg781;
  reg [7:0] y_reg782;
  reg [7:0] y_reg783;
  reg [7:0] y_reg784;
  reg [7:0] y_reg785;
  reg [7:0] y_reg786;
  reg [7:0] y_reg787;
  reg [7:0] y_reg788;
  reg [7:0] y_reg789;
  reg [7:0] y_reg790;
  reg [7:0] y_reg791;
  reg [7:0] y_reg792;
  reg [7:0] y_reg793;
  reg [7:0] y_reg794;
  reg [7:0] y_reg795;
  reg [7:0] y_reg796;
  reg [7:0] y_reg797;
  reg [7:0] y_reg798;
  reg [7:0] y_reg799;
  wire [7:0] t639_b0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t640_b0_G16_mul1_G256_inv0;
  wire [7:0] t641_e0_G256_inv0;
  wire [7:0] t642_p0ls2_G16_inv0_G256_inv0;
  wire [7:0] t643_p0_G16_inv0_G256_inv0;
  wire [7:0] t644_dec_2_inp;
  wire [7:0] t645_q0_G16_inv0_G256_inv0;
  wire [7:0] t646_p0ls1_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t647_q0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t648_dec_3_inp;
  wire [7:0] t649_dec_1_inp;
  wire [7:0] t650_d0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t651_d0_G16_mul1_G256_inv0;
  wire [7:0] t652_b0_G256_inv0;
  wire [7:0] t653_t2;
  wire [7:0] t654_y8_G256_newbasis0;
  wire [7:0] t655_ny8_G256_newbasis0;
  wire [7:0] t656_tempyIntoNegCond8_G256_newbasis0;
  wire [7:0] t657_dec_15_inp;
  wire [7:0] t658_dec_3_inp;
  wire [7:0] t659_dec_1_inp;
  reg [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0_reg117;
  reg [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0_reg118;
  reg [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0_reg119;
  reg [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0_reg120;
  wire [7:0] t608_axorb_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t609_a0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t610_a0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t611_b0_G16_mul1_G256_inv0;
  wire [7:0] t612_e0_G256_inv0;
  wire [7:0] t613_dec_3_inp;
  wire [7:0] t614_dec_2_inp;
  wire [7:0] t615_dec_1_inp;
  wire [7:0] t616_b0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t617_b0_G16_mul1_G256_inv0;
  wire [7:0] t618_e0_G256_inv0;
  wire [7:0] t619_p0ls2_G16_inv0_G256_inv0;
  wire [7:0] t620_q0_G16_inv0_G256_inv0;
  wire [7:0] t621_dec_3_inp;
  wire [7:0] t622_dec_1_inp;
  wire [7:0] t623_cxord_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t624_c0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t625_c0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t626_d0_G16_mul1_G256_inv0;
  wire [7:0] t627_b0_G256_inv0;
  wire [7:0] t628_dec_3_inp;
  wire [7:0] t629_dec_2_inp;
  wire [7:0] t630_dec_1_inp;
  wire [7:0] t631_d0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t632_d0_G16_mul1_G256_inv0;
  wire [7:0] t633_b0_G256_inv0;
  wire [7:0] t634_t2;
  wire [7:0] t635_y8_G256_newbasis0;
  wire [7:0] t636_dec_15_inp;
  wire [7:0] t637_dec_3_inp;
  wire [7:0] t638_dec_1_inp;
  reg [7:0] e0_G4_mul2_G16_mul1_G256_inv0_reg113;
  reg [7:0] e0_G4_mul2_G16_mul1_G256_inv0_reg114;
  reg [7:0] e0_G4_mul2_G16_mul1_G256_inv0_reg115;
  reg [7:0] e0_G4_mul2_G16_mul1_G256_inv0_reg116;
  wire [7:0] t589_a0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t590_a0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t591_b0_G16_mul1_G256_inv0;
  wire [7:0] t592_e0_G256_inv0;
  wire [7:0] t593_p0ls2_G16_inv0_G256_inv0;
  wire [7:0] t594_q0_G16_inv0_G256_inv0;
  wire [7:0] t595_dec_3_inp;
  wire [7:0] t596_dec_2_inp;
  wire [7:0] t597_dec_1_inp;
  wire [7:0] t598_c0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t599_c0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] t600_d0_G16_mul1_G256_inv0;
  wire [7:0] t601_b0_G256_inv0;
  wire [7:0] t602_t2;
  wire [7:0] t603_y8_G256_newbasis0;
  wire [7:0] t604_dec_15_inp;
  wire [7:0] t605_dec_3_inp;
  wire [7:0] t606_dec_2_inp;
  wire [7:0] t607_dec_1_inp;
  reg [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0_reg109;
  reg [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0_reg110;
  reg [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0_reg111;
  reg [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0_reg112;
  wire [7:0] t570_b0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t571_a0_G16_mul1_G256_inv0;
  wire [7:0] t572_a0_0_G16_mul1_G256_inv0;
  wire [7:0] t573_e0_G256_inv0;
  wire [7:0] t574_p0ls2_G16_inv0_G256_inv0;
  wire [7:0] t575_q0_G16_inv0_G256_inv0;
  wire [7:0] t576_dec_12_inp;
  wire [7:0] t577_dec_2_inp;
  wire [7:0] t578_dec_1_inp;
  wire [7:0] t579_d0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t580_c0_G16_mul1_G256_inv0;
  wire [7:0] t581_c0_0_G16_mul1_G256_inv0;
  wire [7:0] t582_b0_G256_inv0;
  wire [7:0] t583_t2;
  wire [7:0] t584_y8_G256_newbasis0;
  wire [7:0] t585_dec_15_inp;
  wire [7:0] t586_dec_12_inp;
  wire [7:0] t587_dec_2_inp;
  wire [7:0] t588_dec_1_inp;
  reg [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0_reg105;
  reg [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0_reg106;
  reg [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0_reg107;
  reg [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0_reg108;
  wire [7:0] t540_axorb_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t541_a0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t542_a0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t543_a0_G16_mul1_G256_inv0;
  wire [7:0] t544_a0_0_G16_mul1_G256_inv0;
  wire [7:0] t545_dec_2_inp;
  wire [7:0] t546_dec_2_inp;
  wire [7:0] t547_dec_1_inp;
  wire [7:0] t548_b0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t549_a0_G16_mul1_G256_inv0;
  wire [7:0] t550_a0_0_G16_mul1_G256_inv0;
  wire [7:0] t551_e0_G256_inv0;
  wire [7:0] t552_dec_12_inp;
  wire [7:0] t553_dec_2_inp;
  wire [7:0] t554_dec_1_inp;
  wire [7:0] t555_cxord_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t556_c0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t557_c0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t558_c0_G16_mul1_G256_inv0;
  wire [7:0] t559_c0_0_G16_mul1_G256_inv0;
  wire [7:0] t560_dec_2_inp;
  wire [7:0] t561_dec_2_inp;
  wire [7:0] t562_dec_1_inp;
  wire [7:0] t563_d0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t564_c0_G16_mul1_G256_inv0;
  wire [7:0] t565_c0_0_G16_mul1_G256_inv0;
  wire [7:0] t566_b0_G256_inv0;
  wire [7:0] t567_dec_12_inp;
  wire [7:0] t568_dec_2_inp;
  wire [7:0] t569_dec_1_inp;
  reg [7:0] e0_G4_mul1_G16_mul1_G256_inv0_reg99;
  reg [7:0] e0_G4_mul1_G16_mul1_G256_inv0_reg100;
  reg [7:0] e0_G4_mul1_G16_mul1_G256_inv0_reg101;
  reg [7:0] e0_G4_mul1_G16_mul1_G256_inv0_reg102;
  reg [7:0] e0_G4_mul1_G16_mul1_G256_inv0_reg103;
  reg [7:0] e0_G4_mul1_G16_mul1_G256_inv0_reg104;
  wire [7:0] t522_a0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t523_a0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t524_a0_G16_mul1_G256_inv0;
  wire [7:0] t525_a0_0_G16_mul1_G256_inv0;
  wire [7:0] t526_e0_G256_inv0;
  wire [7:0] t527_dec_12_inp;
  wire [7:0] t528_dec_2_inp;
  wire [7:0] t529_dec_2_inp;
  wire [7:0] t530_dec_1_inp;
  wire [7:0] t531_c0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t532_c0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] t533_c0_G16_mul1_G256_inv0;
  wire [7:0] t534_c0_0_G16_mul1_G256_inv0;
  wire [7:0] t535_b0_G256_inv0;
  wire [7:0] t536_dec_12_inp;
  wire [7:0] t537_dec_2_inp;
  wire [7:0] t538_dec_2_inp;
  wire [7:0] t539_dec_1_inp;
  reg [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0_reg95;
  reg [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0_reg96;
  reg [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0_reg97;
  reg [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0_reg98;
  wire [7:0] t495_b0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t496_axorb_0_G16_mul1_G256_inv0;
  wire [7:0] t497_a0_G16_mul1_G256_inv0;
  wire [7:0] t498_a0_0_G16_mul1_G256_inv0;
  wire [7:0] t499_e0_G256_inv0;
  wire [7:0] t500_dec_12_inp;
  wire [7:0] t501_dec_2_inp;
  wire [7:0] t502_b0_G16_mul1_G256_inv0;
  wire [7:0] t503_e0_G256_inv0;
  wire [7:0] t504_p0ls2_G16_inv0_G256_inv0;
  wire [7:0] t505_q0_G16_inv0_G256_inv0;
  wire [7:0] t506_dec_3_inp;
  wire [7:0] t507_dec_1_inp;
  wire [7:0] t508_d0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t509_cxord_0_G16_mul1_G256_inv0;
  wire [7:0] t510_c0_G16_mul1_G256_inv0;
  wire [7:0] t511_c0_0_G16_mul1_G256_inv0;
  wire [7:0] t512_b0_G256_inv0;
  wire [7:0] t513_dec_12_inp;
  wire [7:0] t514_dec_2_inp;
  wire [7:0] t515_d0_G16_mul1_G256_inv0;
  wire [7:0] t516_b0_G256_inv0;
  wire [7:0] t517_t2;
  wire [7:0] t518_y8_G256_newbasis0;
  wire [7:0] t519_dec_15_inp;
  wire [7:0] t520_dec_3_inp;
  wire [7:0] t521_dec_1_inp;
  reg [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0_reg91;
  reg [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0_reg92;
  reg [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0_reg93;
  reg [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0_reg94;
  wire [7:0] t461_axorb_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t462_a0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t463_a0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t464_axorb_0_G16_mul1_G256_inv0;
  wire [7:0] t465_a0_G16_mul1_G256_inv0;
  wire [7:0] t466_b0_G16_mul1_G256_inv0;
  wire [7:0] t467_dec_2_inp;
  wire [7:0] t468_dec_1_inp;
  wire [7:0] t469_b0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t470_axorb_0_G16_mul1_G256_inv0;
  wire [7:0] t471_a0_G16_mul1_G256_inv0;
  wire [7:0] t472_a0_0_G16_mul1_G256_inv0;
  wire [7:0] t473_dec_2_inp;
  wire [7:0] t474_b0_G16_mul1_G256_inv0;
  wire [7:0] t475_e0_G256_inv0;
  wire [7:0] t476_dec_3_inp;
  wire [7:0] t477_dec_1_inp;
  wire [7:0] t478_cxord_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t479_c0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t480_c0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t481_cxord_0_G16_mul1_G256_inv0;
  wire [7:0] t482_c0_G16_mul1_G256_inv0;
  wire [7:0] t483_d0_G16_mul1_G256_inv0;
  wire [7:0] t484_dec_2_inp;
  wire [7:0] t485_dec_1_inp;
  wire [7:0] t486_d0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t487_cxord_0_G16_mul1_G256_inv0;
  wire [7:0] t488_c0_G16_mul1_G256_inv0;
  wire [7:0] t489_c0_0_G16_mul1_G256_inv0;
  wire [7:0] t490_dec_2_inp;
  wire [7:0] t491_d0_G16_mul1_G256_inv0;
  wire [7:0] t492_b0_G256_inv0;
  wire [7:0] t493_dec_3_inp;
  wire [7:0] t494_dec_1_inp;
  reg [7:0] e0_G4_mul0_G16_mul1_G256_inv0_reg85;
  reg [7:0] e0_G4_mul0_G16_mul1_G256_inv0_reg86;
  reg [7:0] e0_G4_mul0_G16_mul1_G256_inv0_reg87;
  reg [7:0] e0_G4_mul0_G16_mul1_G256_inv0_reg88;
  reg [7:0] e0_G4_mul0_G16_mul1_G256_inv0_reg89;
  reg [7:0] e0_G4_mul0_G16_mul1_G256_inv0_reg90;
  wire [7:0] t439_a0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t440_a0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t441_axorb_0_G16_mul1_G256_inv0;
  wire [7:0] t442_a0_G16_mul1_G256_inv0;
  wire [7:0] t443_a0_0_G16_mul1_G256_inv0;
  wire [7:0] t444_dec_2_inp;
  wire [7:0] t445_b0_G16_mul1_G256_inv0;
  wire [7:0] t446_e0_G256_inv0;
  wire [7:0] t447_dec_3_inp;
  wire [7:0] t448_dec_2_inp;
  wire [7:0] t449_dec_1_inp;
  wire [7:0] t450_c0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t451_c0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] t452_cxord_0_G16_mul1_G256_inv0;
  wire [7:0] t453_c0_G16_mul1_G256_inv0;
  wire [7:0] t454_c0_0_G16_mul1_G256_inv0;
  wire [7:0] t455_dec_2_inp;
  wire [7:0] t456_d0_G16_mul1_G256_inv0;
  wire [7:0] t457_b0_G256_inv0;
  wire [7:0] t458_dec_3_inp;
  wire [7:0] t459_dec_2_inp;
  wire [7:0] t460_dec_1_inp;
  reg [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0_reg81;
  reg [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0_reg82;
  reg [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0_reg83;
  reg [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0_reg84;
  wire [7:0] t417_b0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t418_e0_G16_inv0_G256_inv0;
  wire [7:0] t419_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t420_b0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t421_c0xord0_G16_inv0_G256_inv0;
  wire [7:0] t422_dec_1_inp;
  wire [7:0] t423_dec_1_inp;
  wire [7:0] t424_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t425_a0_0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t426_c0xord0_G16_inv0_G256_inv0;
  wire [7:0] t427_dec_2_inp;
  wire [7:0] t428_dec_1_inp;
  wire [7:0] t429_dec_1_inp;
  wire [7:0] t430_d0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t431_a0_G16_inv0_G256_inv0;
  wire [7:0] t432_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t433_c0xord0_G256_inv0;
  wire [7:0] t434_c0_G256_inv0;
  wire [7:0] t435_d0_G256_inv0;
  wire [7:0] t436_dec_12_inp;
  wire [7:0] t437_dec_2_inp;
  wire [7:0] t438_dec_1_inp;
  reg [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0_reg77;
  reg [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0_reg78;
  reg [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0_reg79;
  reg [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0_reg80;
  wire [7:0] t385_axorb_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t386_a0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t387_a0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t388_e0_G16_inv0_G256_inv0;
  wire [7:0] t389_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t390_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t391_dec_2_inp;
  wire [7:0] t392_dec_1_inp;
  wire [7:0] t393_b0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t394_e0_G16_inv0_G256_inv0;
  wire [7:0] t395_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t396_b0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t397_dec_1_inp;
  wire [7:0] t398_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t399_a0_0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t400_dec_1_inp;
  wire [7:0] t401_dec_1_inp;
  wire [7:0] t402_cxord_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t403_c0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t404_c0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t405_a0_G16_inv0_G256_inv0;
  wire [7:0] t406_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t407_dec_2_inp;
  wire [7:0] t408_dec_2_inp;
  wire [7:0] t409_dec_1_inp;
  wire [7:0] t410_d0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t411_a0_G16_inv0_G256_inv0;
  wire [7:0] t412_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t413_c0xord0_G256_inv0;
  wire [7:0] t414_dec_12_inp;
  wire [7:0] t415_dec_2_inp;
  wire [7:0] t416_dec_1_inp;
  reg [7:0] e0_G4_mul5_G16_inv0_G256_inv0_reg71;
  reg [7:0] e0_G4_mul5_G16_inv0_G256_inv0_reg72;
  reg [7:0] e0_G4_mul5_G16_inv0_G256_inv0_reg73;
  reg [7:0] e0_G4_mul5_G16_inv0_G256_inv0_reg74;
  reg [7:0] e0_G4_mul5_G16_inv0_G256_inv0_reg75;
  reg [7:0] e0_G4_mul5_G16_inv0_G256_inv0_reg76;
  wire [7:0] t365_a0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t366_a0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t367_e0_G16_inv0_G256_inv0;
  wire [7:0] t368_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t369_b0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t370_dec_1_inp;
  wire [7:0] t371_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t372_a0_0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t373_dec_1_inp;
  wire [7:0] t374_dec_2_inp;
  wire [7:0] t375_dec_1_inp;
  wire [7:0] t376_c0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t377_c0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] t378_a0_G16_inv0_G256_inv0;
  wire [7:0] t379_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t380_c0xord0_G256_inv0;
  wire [7:0] t381_dec_12_inp;
  wire [7:0] t382_dec_2_inp;
  wire [7:0] t383_dec_2_inp;
  wire [7:0] t384_dec_1_inp;
  reg [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0_reg67;
  reg [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0_reg68;
  reg [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0_reg69;
  reg [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0_reg70;
  wire [7:0] t341_b0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t342_e0_G16_inv0_G256_inv0;
  wire [7:0] t343_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t344_b0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t345_c0xord0_G16_inv0_G256_inv0;
  wire [7:0] t346_dec_1_inp;
  wire [7:0] t347_dec_1_inp;
  wire [7:0] t348_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t349_a0_0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t350_c0xord0_G16_inv0_G256_inv0;
  wire [7:0] t351_dec_2_inp;
  wire [7:0] t352_dec_1_inp;
  wire [7:0] t353_dec_1_inp;
  wire [7:0] t354_d0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t355_b0_G16_inv0_G256_inv0;
  wire [7:0] t356_c0xord0_G256_inv0;
  wire [7:0] t357_c0_G256_inv0;
  wire [7:0] t358_p0ls2_G16_sq_scl0_G256_inv0;
  wire [7:0] t359_q0_G16_sq_scl0_G256_inv0;
  wire [7:0] t360_d0_G256_inv0;
  wire [7:0] t361_p0ls2_G16_mul0_G256_inv0;
  wire [7:0] t362_q0_G16_mul0_G256_inv0;
  wire [7:0] t363_dec_3_inp;
  wire [7:0] t364_dec_1_inp;
  reg [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0_reg63;
  reg [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0_reg64;
  reg [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0_reg65;
  reg [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0_reg66;
  wire [7:0] t309_axorb_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t310_a0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t311_a0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t312_e0_G16_inv0_G256_inv0;
  wire [7:0] t313_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t314_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t315_dec_2_inp;
  wire [7:0] t316_dec_1_inp;
  wire [7:0] t317_b0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t318_e0_G16_inv0_G256_inv0;
  wire [7:0] t319_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t320_b0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t321_dec_1_inp;
  wire [7:0] t322_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t323_a0_0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t324_dec_1_inp;
  wire [7:0] t325_dec_1_inp;
  wire [7:0] t326_cxord_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t327_c0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t328_c0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t329_b0_G16_inv0_G256_inv0;
  wire [7:0] t330_c0xord0_G256_inv0;
  wire [7:0] t331_dec_3_inp;
  wire [7:0] t332_dec_2_inp;
  wire [7:0] t333_dec_1_inp;
  wire [7:0] t334_d0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t335_b0_G16_inv0_G256_inv0;
  wire [7:0] t336_c0xord0_G256_inv0;
  wire [7:0] t337_c0_G256_inv0;
  wire [7:0] t338_d0_G256_inv0;
  wire [7:0] t339_dec_3_inp;
  wire [7:0] t340_dec_1_inp;
  reg [7:0] e0_G4_mul4_G16_inv0_G256_inv0_reg59;
  reg [7:0] e0_G4_mul4_G16_inv0_G256_inv0_reg60;
  reg [7:0] e0_G4_mul4_G16_inv0_G256_inv0_reg61;
  reg [7:0] e0_G4_mul4_G16_inv0_G256_inv0_reg62;
  wire [7:0] t289_a0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t290_a0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t291_e0_G16_inv0_G256_inv0;
  wire [7:0] t292_b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t293_b0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t294_dec_1_inp;
  wire [7:0] t295_a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t296_a0_0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] t297_dec_1_inp;
  wire [7:0] t298_dec_2_inp;
  wire [7:0] t299_dec_1_inp;
  wire [7:0] t300_c0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t301_c0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] t302_b0_G16_inv0_G256_inv0;
  wire [7:0] t303_c0xord0_G256_inv0;
  wire [7:0] t304_c0_G256_inv0;
  wire [7:0] t305_d0_G256_inv0;
  wire [7:0] t306_dec_3_inp;
  wire [7:0] t307_dec_2_inp;
  wire [7:0] t308_dec_1_inp;
  reg [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0_reg55;
  reg [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0_reg56;
  reg [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0_reg57;
  reg [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0_reg58;
  wire [7:0] t269_b0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t270_a0_G16_inv0_G256_inv0;
  wire [7:0] t271_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t272_c0xord0_G256_inv0;
  wire [7:0] t273_c0_G256_inv0;
  wire [7:0] t274_d0_G256_inv0;
  wire [7:0] t275_dec_12_inp;
  wire [7:0] t276_dec_2_inp;
  wire [7:0] t277_dec_1_inp;
  wire [7:0] t278_d0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t279_b0_G16_inv0_G256_inv0;
  wire [7:0] t280_c0xord0_G256_inv0;
  wire [7:0] t281_c0_G256_inv0;
  wire [7:0] t282_p0ls2_G16_sq_scl0_G256_inv0;
  wire [7:0] t283_q0_G16_sq_scl0_G256_inv0;
  wire [7:0] t284_d0_G256_inv0;
  wire [7:0] t285_p0ls2_G16_mul0_G256_inv0;
  wire [7:0] t286_q0_G16_mul0_G256_inv0;
  wire [7:0] t287_dec_3_inp;
  wire [7:0] t288_dec_1_inp;
  reg [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0_reg51;
  reg [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0_reg52;
  reg [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0_reg53;
  reg [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0_reg54;
  wire [7:0] t239_axorb_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t240_a0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t241_a0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t242_a0_G16_inv0_G256_inv0;
  wire [7:0] t243_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t244_dec_2_inp;
  wire [7:0] t245_dec_2_inp;
  wire [7:0] t246_dec_1_inp;
  wire [7:0] t247_b0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t248_a0_G16_inv0_G256_inv0;
  wire [7:0] t249_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t250_c0xord0_G256_inv0;
  wire [7:0] t251_dec_12_inp;
  wire [7:0] t252_dec_2_inp;
  wire [7:0] t253_dec_1_inp;
  wire [7:0] t254_cxord_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t255_c0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t256_c0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t257_b0_G16_inv0_G256_inv0;
  wire [7:0] t258_c0xord0_G256_inv0;
  wire [7:0] t259_dec_3_inp;
  wire [7:0] t260_dec_2_inp;
  wire [7:0] t261_dec_1_inp;
  wire [7:0] t262_d0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t263_b0_G16_inv0_G256_inv0;
  wire [7:0] t264_c0xord0_G256_inv0;
  wire [7:0] t265_c0_G256_inv0;
  wire [7:0] t266_d0_G256_inv0;
  wire [7:0] t267_dec_3_inp;
  wire [7:0] t268_dec_1_inp;
  reg [7:0] e0_G4_mul3_G16_inv0_G256_inv0_reg45;
  reg [7:0] e0_G4_mul3_G16_inv0_G256_inv0_reg46;
  reg [7:0] e0_G4_mul3_G16_inv0_G256_inv0_reg47;
  reg [7:0] e0_G4_mul3_G16_inv0_G256_inv0_reg48;
  reg [7:0] e0_G4_mul3_G16_inv0_G256_inv0_reg49;
  reg [7:0] e0_G4_mul3_G16_inv0_G256_inv0_reg50;
  wire [7:0] t221_a0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t222_a0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t223_a0_G16_inv0_G256_inv0;
  wire [7:0] t224_a0_0_G16_inv0_G256_inv0;
  wire [7:0] t225_c0xord0_G256_inv0;
  wire [7:0] t226_dec_12_inp;
  wire [7:0] t227_dec_2_inp;
  wire [7:0] t228_dec_2_inp;
  wire [7:0] t229_dec_1_inp;
  wire [7:0] t230_c0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t231_c0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] t232_b0_G16_inv0_G256_inv0;
  wire [7:0] t233_c0xord0_G256_inv0;
  wire [7:0] t234_c0_G256_inv0;
  wire [7:0] t235_d0_G256_inv0;
  wire [7:0] t236_dec_3_inp;
  wire [7:0] t237_dec_2_inp;
  wire [7:0] t238_dec_1_inp;
  reg [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0_reg41;
  reg [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0_reg42;
  reg [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0_reg43;
  reg [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0_reg44;
  wire [7:0] t201_b0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t202_b0_G16_mul0_G256_inv0;
  wire [7:0] t203_a0_G256_inv0;
  wire [7:0] t204_a0_0_G256_inv0;
  wire [7:0] t205_t2;
  wire [7:0] t206_y8_G256_newbasis0;
  wire [7:0] t207_dec_240_inp;
  wire [7:0] t208_dec_4_inp;
  wire [7:0] t209_dec_3_inp;
  wire [7:0] t210_dec_1_inp;
  wire [7:0] t211_d0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t212_d0_G16_mul0_G256_inv0;
  wire [7:0] t213_b0_G256_inv0;
  wire [7:0] t214_t2;
  wire [7:0] t215_y8_G256_newbasis0;
  wire [7:0] t216_ny8_G256_newbasis0;
  wire [7:0] t217_tempyIntoNegCond8_G256_newbasis0;
  wire [7:0] t218_dec_15_inp;
  wire [7:0] t219_dec_3_inp;
  wire [7:0] t220_dec_1_inp;
  reg [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0_reg37;
  reg [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0_reg38;
  reg [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0_reg39;
  reg [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0_reg40;
  wire [7:0] t170_axorb_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t171_a0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t172_a0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t173_b0_G16_mul0_G256_inv0;
  wire [7:0] t174_a0_G256_inv0;
  wire [7:0] t175_dec_3_inp;
  wire [7:0] t176_dec_2_inp;
  wire [7:0] t177_dec_1_inp;
  wire [7:0] t178_b0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t179_b0_G16_mul0_G256_inv0;
  wire [7:0] t180_a0_G256_inv0;
  wire [7:0] t181_a0_0_G256_inv0;
  wire [7:0] t182_dec_4_inp;
  wire [7:0] t183_dec_3_inp;
  wire [7:0] t184_dec_1_inp;
  wire [7:0] t185_cxord_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t186_c0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t187_c0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t188_d0_G16_mul0_G256_inv0;
  wire [7:0] t189_b0_G256_inv0;
  wire [7:0] t190_dec_3_inp;
  wire [7:0] t191_dec_2_inp;
  wire [7:0] t192_dec_1_inp;
  wire [7:0] t193_d0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t194_d0_G16_mul0_G256_inv0;
  wire [7:0] t195_b0_G256_inv0;
  wire [7:0] t196_t2;
  wire [7:0] t197_y8_G256_newbasis0;
  wire [7:0] t198_dec_15_inp;
  wire [7:0] t199_dec_3_inp;
  wire [7:0] t200_dec_1_inp;
  reg [7:0] e0_G4_mul2_G16_mul0_G256_inv0_reg31;
  reg [7:0] e0_G4_mul2_G16_mul0_G256_inv0_reg32;
  reg [7:0] e0_G4_mul2_G16_mul0_G256_inv0_reg33;
  reg [7:0] e0_G4_mul2_G16_mul0_G256_inv0_reg34;
  reg [7:0] e0_G4_mul2_G16_mul0_G256_inv0_reg35;
  reg [7:0] e0_G4_mul2_G16_mul0_G256_inv0_reg36;
  wire [7:0] t151_a0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t152_a0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t153_b0_G16_mul0_G256_inv0;
  wire [7:0] t154_a0_G256_inv0;
  wire [7:0] t155_a0_0_G256_inv0;
  wire [7:0] t156_dec_4_inp;
  wire [7:0] t157_dec_3_inp;
  wire [7:0] t158_dec_2_inp;
  wire [7:0] t159_dec_1_inp;
  wire [7:0] t160_c0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t161_c0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] t162_d0_G16_mul0_G256_inv0;
  wire [7:0] t163_b0_G256_inv0;
  wire [7:0] t164_t2;
  wire [7:0] t165_y8_G256_newbasis0;
  wire [7:0] t166_dec_15_inp;
  wire [7:0] t167_dec_3_inp;
  wire [7:0] t168_dec_2_inp;
  wire [7:0] t169_dec_1_inp;
  reg [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0_reg27;
  reg [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0_reg28;
  reg [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0_reg29;
  reg [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0_reg30;
  wire [7:0] t132_b0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t133_a0_G16_mul0_G256_inv0;
  wire [7:0] t134_a0_0_G16_mul0_G256_inv0;
  wire [7:0] t135_a0_G256_inv0;
  wire [7:0] t136_a0_0_G256_inv0;
  wire [7:0] t137_dec_4_inp;
  wire [7:0] t138_dec_12_inp;
  wire [7:0] t139_dec_2_inp;
  wire [7:0] t140_dec_1_inp;
  wire [7:0] t141_d0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t142_c0_G16_mul0_G256_inv0;
  wire [7:0] t143_c0_0_G16_mul0_G256_inv0;
  wire [7:0] t144_b0_G256_inv0;
  wire [7:0] t145_t2;
  wire [7:0] t146_y8_G256_newbasis0;
  wire [7:0] t147_dec_15_inp;
  wire [7:0] t148_dec_12_inp;
  wire [7:0] t149_dec_2_inp;
  wire [7:0] t150_dec_1_inp;
  reg [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0_reg23;
  reg [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0_reg24;
  reg [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0_reg25;
  reg [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0_reg26;
  wire [7:0] t102_axorb_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t103_a0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t104_a0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t105_a0_G16_mul0_G256_inv0;
  wire [7:0] t106_a0_0_G16_mul0_G256_inv0;
  wire [7:0] t107_dec_2_inp;
  wire [7:0] t108_dec_2_inp;
  wire [7:0] t109_dec_1_inp;
  wire [7:0] t110_b0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t111_a0_G16_mul0_G256_inv0;
  wire [7:0] t112_a0_0_G16_mul0_G256_inv0;
  wire [7:0] t113_a0_G256_inv0;
  wire [7:0] t114_dec_12_inp;
  wire [7:0] t115_dec_2_inp;
  wire [7:0] t116_dec_1_inp;
  wire [7:0] t117_cxord_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t118_c0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t119_c0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t120_c0_G16_mul0_G256_inv0;
  wire [7:0] t121_c0_0_G16_mul0_G256_inv0;
  wire [7:0] t122_dec_2_inp;
  wire [7:0] t123_dec_2_inp;
  wire [7:0] t124_dec_1_inp;
  wire [7:0] t125_d0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t126_c0_G16_mul0_G256_inv0;
  wire [7:0] t127_c0_0_G16_mul0_G256_inv0;
  wire [7:0] t128_b0_G256_inv0;
  wire [7:0] t129_dec_12_inp;
  wire [7:0] t130_dec_2_inp;
  wire [7:0] t131_dec_1_inp;
  reg [7:0] e0_G4_mul1_G16_mul0_G256_inv0_reg17;
  reg [7:0] e0_G4_mul1_G16_mul0_G256_inv0_reg18;
  reg [7:0] e0_G4_mul1_G16_mul0_G256_inv0_reg19;
  reg [7:0] e0_G4_mul1_G16_mul0_G256_inv0_reg20;
  reg [7:0] e0_G4_mul1_G16_mul0_G256_inv0_reg21;
  reg [7:0] e0_G4_mul1_G16_mul0_G256_inv0_reg22;
  wire [7:0] t84_a0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t85_a0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t86_a0_G16_mul0_G256_inv0;
  wire [7:0] t87_a0_0_G16_mul0_G256_inv0;
  wire [7:0] t88_a0_G256_inv0;
  wire [7:0] t89_dec_12_inp;
  wire [7:0] t90_dec_2_inp;
  wire [7:0] t91_dec_2_inp;
  wire [7:0] t92_dec_1_inp;
  wire [7:0] t93_c0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t94_c0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] t95_c0_G16_mul0_G256_inv0;
  wire [7:0] t96_c0_0_G16_mul0_G256_inv0;
  wire [7:0] t97_b0_G256_inv0;
  wire [7:0] t98_dec_12_inp;
  wire [7:0] t99_dec_2_inp;
  wire [7:0] t100_dec_2_inp;
  wire [7:0] t101_dec_1_inp;
  reg [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0_reg13;
  reg [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0_reg14;
  reg [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0_reg15;
  reg [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0_reg16;
  wire [7:0] t57_b0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t58_axorb_0_G16_mul0_G256_inv0;
  wire [7:0] t59_a0_G16_mul0_G256_inv0;
  wire [7:0] t60_a0_0_G16_mul0_G256_inv0;
  wire [7:0] t61_a0_G256_inv0;
  wire [7:0] t62_dec_12_inp;
  wire [7:0] t63_dec_2_inp;
  wire [7:0] t64_b0_G16_mul0_G256_inv0;
  wire [7:0] t65_a0_G256_inv0;
  wire [7:0] t66_a0_0_G256_inv0;
  wire [7:0] t67_dec_4_inp;
  wire [7:0] t68_dec_3_inp;
  wire [7:0] t69_dec_1_inp;
  wire [7:0] t70_d0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t71_cxord_0_G16_mul0_G256_inv0;
  wire [7:0] t72_c0_G16_mul0_G256_inv0;
  wire [7:0] t73_c0_0_G16_mul0_G256_inv0;
  wire [7:0] t74_b0_G256_inv0;
  wire [7:0] t75_dec_12_inp;
  wire [7:0] t76_dec_2_inp;
  wire [7:0] t77_d0_G16_mul0_G256_inv0;
  wire [7:0] t78_b0_G256_inv0;
  wire [7:0] t79_t2;
  wire [7:0] t80_y8_G256_newbasis0;
  wire [7:0] t81_dec_15_inp;
  wire [7:0] t82_dec_3_inp;
  wire [7:0] t83_dec_1_inp;
  reg [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0_reg9;
  reg [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0_reg10;
  reg [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0_reg11;
  reg [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0_reg12;
  wire [7:0] t23_axorb_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t24_a0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t25_a0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t26_axorb_0_G16_mul0_G256_inv0;
  wire [7:0] t27_a0_G16_mul0_G256_inv0;
  wire [7:0] t28_b0_G16_mul0_G256_inv0;
  wire [7:0] t29_dec_2_inp;
  wire [7:0] t30_dec_1_inp;
  wire [7:0] t31_b0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t32_axorb_0_G16_mul0_G256_inv0;
  wire [7:0] t33_a0_G16_mul0_G256_inv0;
  wire [7:0] t34_a0_0_G16_mul0_G256_inv0;
  wire [7:0] t35_dec_2_inp;
  wire [7:0] t36_b0_G16_mul0_G256_inv0;
  wire [7:0] t37_a0_G256_inv0;
  wire [7:0] t38_dec_3_inp;
  wire [7:0] t39_dec_1_inp;
  wire [7:0] t40_cxord_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t41_c0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t42_c0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t43_cxord_0_G16_mul0_G256_inv0;
  wire [7:0] t44_c0_G16_mul0_G256_inv0;
  wire [7:0] t45_d0_G16_mul0_G256_inv0;
  wire [7:0] t46_dec_2_inp;
  wire [7:0] t47_dec_1_inp;
  wire [7:0] t48_d0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t49_cxord_0_G16_mul0_G256_inv0;
  wire [7:0] t50_c0_G16_mul0_G256_inv0;
  wire [7:0] t51_c0_0_G16_mul0_G256_inv0;
  wire [7:0] t52_dec_2_inp;
  wire [7:0] t53_d0_G16_mul0_G256_inv0;
  wire [7:0] t54_b0_G256_inv0;
  wire [7:0] t55_dec_3_inp;
  wire [7:0] t56_dec_1_inp;
  reg [7:0] e0_G4_mul0_G16_mul0_G256_inv0_reg5;
  reg [7:0] e0_G4_mul0_G16_mul0_G256_inv0_reg6;
  reg [7:0] e0_G4_mul0_G16_mul0_G256_inv0_reg7;
  reg [7:0] e0_G4_mul0_G16_mul0_G256_inv0_reg8;
  wire [7:0] t1_a0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t2_a0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t3_axorb_0_G16_mul0_G256_inv0;
  wire [7:0] t4_a0_G16_mul0_G256_inv0;
  wire [7:0] t5_a0_0_G16_mul0_G256_inv0;
  wire [7:0] t6_dec_2_inp;
  wire [7:0] t7_b0_G16_mul0_G256_inv0;
  wire [7:0] t8_a0_G256_inv0;
  wire [7:0] t9_dec_3_inp;
  wire [7:0] t10_dec_2_inp;
  wire [7:0] t11_dec_1_inp;
  wire [7:0] t12_c0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t13_c0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] t14_cxord_0_G16_mul0_G256_inv0;
  wire [7:0] t15_c0_G16_mul0_G256_inv0;
  wire [7:0] t16_c0_0_G16_mul0_G256_inv0;
  wire [7:0] t17_dec_2_inp;
  wire [7:0] t18_d0_G16_mul0_G256_inv0;
  wire [7:0] t19_b0_G256_inv0;
  wire [7:0] t20_dec_3_inp;
  wire [7:0] t21_dec_2_inp;
  wire [7:0] t22_dec_1_inp;
  reg [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0_reg1;
  reg [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0_reg2;
  reg [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0_reg3;
  reg [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0_reg4;
  input clk;
  input [7:0] t;
  input [7:0] dec_0;
  input [7:0] dec_1;
  input [7:0] dec_255;
  input [7:0] dec_169;
  input [7:0] dec_129;
  input [7:0] dec_9;
  input [7:0] dec_72;
  input [7:0] dec_242;
  input [7:0] dec_243;
  input [7:0] dec_152;
  input [7:0] dec_240;
  input [7:0] dec_4;
  input [7:0] dec_15;
  input [7:0] dec_12;
  input [7:0] dec_2;
  input [7:0] dec_3;
  input [7:0] dec_36;
  input [7:0] dec_220;
  input [7:0] dec_11;
  input [7:0] dec_158;
  input [7:0] dec_45;
  input [7:0] dec_88;
  input [7:0] dec_99;
  input [20:0] r;
  output [7:0] y;reg [7:0] y;
  wire [7:0] dec_99_inp;
  wire [7:0] dec_88_inp;
  wire [7:0] dec_45_inp;
  wire [7:0] dec_158_inp;
  wire [7:0] dec_11_inp;
  wire [7:0] dec_220_inp;
  wire [7:0] dec_36_inp;
  wire [7:0] dec_3_inp;
  wire [7:0] dec_2_inp;
  wire [7:0] dec_12_inp;
  wire [7:0] dec_15_inp;
  wire [7:0] dec_4_inp;
  wire [7:0] dec_240_inp;
  wire [7:0] dec_152_inp;
  wire [7:0] dec_243_inp;
  wire [7:0] dec_242_inp;
  wire [7:0] dec_72_inp;
  wire [7:0] dec_9_inp;
  wire [7:0] dec_129_inp;
  wire [7:0] dec_169_inp;
  wire [7:0] dec_255_inp;
  wire [7:0] dec_1_inp;
  wire [7:0] dec_0_inp;
  wire [7:0] t_inp;
  wire [7:0] y_G256_newbasis0;
  wire [7:0] tempy1_G256_newbasis0;
  wire [7:0] cond1_G256_newbasis0;
  wire [7:0] negCond1_G256_newbasis0;
  wire [7:0] yxorb1_G256_newbasis0;
  wire [7:0] ny1_G256_newbasis0;
  wire [7:0] tempyIntoNegCond1_G256_newbasis0;
  wire [7:0] y1_G256_newbasis0;
  wire [7:0] x1_G256_newbasis0;
  wire [7:0] tempy2_G256_newbasis0;
  wire [7:0] cond2_G256_newbasis0;
  wire [7:0] negCond2_G256_newbasis0;
  wire [7:0] yxorb2_G256_newbasis0;
  wire [7:0] ny2_G256_newbasis0;
  wire [7:0] tempyIntoNegCond2_G256_newbasis0;
  wire [7:0] y2_G256_newbasis0;
  wire [7:0] x2_G256_newbasis0;
  wire [7:0] tempy3_G256_newbasis0;
  wire [7:0] cond3_G256_newbasis0;
  wire [7:0] negCond3_G256_newbasis0;
  wire [7:0] yxorb3_G256_newbasis0;
  wire [7:0] ny3_G256_newbasis0;
  wire [7:0] tempyIntoNegCond3_G256_newbasis0;
  wire [7:0] y3_G256_newbasis0;
  wire [7:0] x3_G256_newbasis0;
  wire [7:0] tempy4_G256_newbasis0;
  wire [7:0] cond4_G256_newbasis0;
  wire [7:0] negCond4_G256_newbasis0;
  wire [7:0] yxorb4_G256_newbasis0;
  wire [7:0] ny4_G256_newbasis0;
  wire [7:0] tempyIntoNegCond4_G256_newbasis0;
  wire [7:0] y4_G256_newbasis0;
  wire [7:0] x4_G256_newbasis0;
  wire [7:0] tempy5_G256_newbasis0;
  wire [7:0] cond5_G256_newbasis0;
  wire [7:0] negCond5_G256_newbasis0;
  wire [7:0] yxorb5_G256_newbasis0;
  wire [7:0] ny5_G256_newbasis0;
  wire [7:0] tempyIntoNegCond5_G256_newbasis0;
  wire [7:0] y5_G256_newbasis0;
  wire [7:0] x5_G256_newbasis0;
  wire [7:0] tempy6_G256_newbasis0;
  wire [7:0] cond6_G256_newbasis0;
  wire [7:0] negCond6_G256_newbasis0;
  wire [7:0] yxorb6_G256_newbasis0;
  wire [7:0] ny6_G256_newbasis0;
  wire [7:0] tempyIntoNegCond6_G256_newbasis0;
  wire [7:0] y6_G256_newbasis0;
  wire [7:0] x6_G256_newbasis0;
  wire [7:0] tempy7_G256_newbasis0;
  wire [7:0] cond7_G256_newbasis0;
  wire [7:0] negCond7_G256_newbasis0;
  wire [7:0] yxorb7_G256_newbasis0;
  wire [7:0] ny7_G256_newbasis0;
  wire [7:0] tempyIntoNegCond7_G256_newbasis0;
  wire [7:0] y7_G256_newbasis0;
  wire [7:0] x7_G256_newbasis0;
  wire [7:0] tempy8_G256_newbasis0;
  wire [7:0] cond8_G256_newbasis0;
  wire [7:0] negCond8_G256_newbasis0;
  wire [7:0] yxorb8_G256_newbasis0;
  wire [7:0] ny8_G256_newbasis0;
  wire [7:0] tempyIntoNegCond8_G256_newbasis0;
  wire [7:0] y8_G256_newbasis0;
  wire [7:0] x8_G256_newbasis0;
  wire [7:0] t2;
  wire [7:0] a0_0_G256_inv0;
  wire [7:0] a0_G256_inv0;
  wire [7:0] b0_G256_inv0;
  wire [7:0] a0xorb0_G256_inv0;
  wire [7:0] a0_0_G16_sq_scl0_G256_inv0;
  wire [7:0] a0_G16_sq_scl0_G256_inv0;
  wire [7:0] b0_G16_sq_scl0_G256_inv0;
  wire [7:0] p0_0_G16_sq_scl0_G256_inv0;
  wire [7:0] a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
  wire [7:0] a0_G4_sq0_G16_sq_scl0_G256_inv0;
  wire [7:0] b0_G4_sq0_G16_sq_scl0_G256_inv0;
  wire [7:0] b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
  wire [7:0] p0_G16_sq_scl0_G256_inv0;
  wire [7:0] a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
  wire [7:0] a0_G4_sq1_G16_sq_scl0_G256_inv0;
  wire [7:0] b0_G4_sq1_G16_sq_scl0_G256_inv0;
  wire [7:0] b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
  wire [7:0] q0_0_G16_sq_scl0_G256_inv0;
  wire [7:0] a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  wire [7:0] a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  wire [7:0] b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  wire [7:0] p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  wire [7:0] q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  wire [7:0] p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
  wire [7:0] q0_G16_sq_scl0_G256_inv0;
  wire [7:0] p0ls2_G16_sq_scl0_G256_inv0;
  wire [7:0] c0_G256_inv0;
  wire [7:0] a0_0_G16_mul0_G256_inv0;
  wire [7:0] a0_G16_mul0_G256_inv0;
  wire [7:0] b0_G16_mul0_G256_inv0;
  wire [7:0] c0_0_G16_mul0_G256_inv0;
  wire [7:0] c0_G16_mul0_G256_inv0;
  wire [7:0] d0_G16_mul0_G256_inv0;
  wire [7:0] axorb_0_G16_mul0_G256_inv0;
  wire [7:0] cxord_0_G16_mul0_G256_inv0;
  wire [7:0] a0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] a0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] b0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] c0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] c0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] d0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] axorb_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] cxord_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] e0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] p0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] q0_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] p0ls1_G4_mul0_G16_mul0_G256_inv0;
  wire [7:0] e0_G16_mul0_G256_inv0;
  wire [7:0] a0_0_G4_scl_N0_G16_mul0_G256_inv0;
  wire [7:0] a0_G4_scl_N0_G16_mul0_G256_inv0;
  wire [7:0] b0_G4_scl_N0_G16_mul0_G256_inv0;
  wire [7:0] p0_G4_scl_N0_G16_mul0_G256_inv0;
  wire [7:0] q0_G4_scl_N0_G16_mul0_G256_inv0;
  wire [7:0] p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
  wire [7:0] e01_G16_mul0_G256_inv0;
  wire [7:0] a0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] a0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] b0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] c0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] c0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] d0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] axorb_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] cxord_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] e0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] p0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] q0_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] p0ls1_G4_mul1_G16_mul0_G256_inv0;
  wire [7:0] p0_0_G16_mul0_G256_inv0;
  wire [7:0] p0_G16_mul0_G256_inv0;
  wire [7:0] a0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] a0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] b0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] c0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] c0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] d0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] axorb_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] cxord_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] e0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] p0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] q0_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] p0ls1_G4_mul2_G16_mul0_G256_inv0;
  wire [7:0] q0_0_G16_mul0_G256_inv0;
  wire [7:0] q0_G16_mul0_G256_inv0;
  wire [7:0] p0ls2_G16_mul0_G256_inv0;
  wire [7:0] d0_G256_inv0;
  wire [7:0] c0xord0_G256_inv0;
  wire [7:0] a0_0_G16_inv0_G256_inv0;
  wire [7:0] a0_G16_inv0_G256_inv0;
  wire [7:0] b0_G16_inv0_G256_inv0;
  wire [7:0] a0xorb0_G16_inv0_G256_inv0;
  wire [7:0] a0_0_G4_sq2_G16_inv0_G256_inv0;
  wire [7:0] a0_G4_sq2_G16_inv0_G256_inv0;
  wire [7:0] b0_G4_sq2_G16_inv0_G256_inv0;
  wire [7:0] b0ls1_G4_sq2_G16_inv0_G256_inv0;
  wire [7:0] c0_0_G16_inv0_G256_inv0;
  wire [7:0] a0_0_G4_scl_N1_G16_inv0_G256_inv0;
  wire [7:0] a0_G4_scl_N1_G16_inv0_G256_inv0;
  wire [7:0] b0_G4_scl_N1_G16_inv0_G256_inv0;
  wire [7:0] p0_G4_scl_N1_G16_inv0_G256_inv0;
  wire [7:0] q0_G4_scl_N1_G16_inv0_G256_inv0;
  wire [7:0] p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
  wire [7:0] c0_G16_inv0_G256_inv0;
  wire [7:0] a0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] a0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] b0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] c0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] c0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] d0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] axorb_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] cxord_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] e0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] p0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] q0_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] p0ls1_G4_mul3_G16_inv0_G256_inv0;
  wire [7:0] d0_G16_inv0_G256_inv0;
  wire [7:0] c0xord0_G16_inv0_G256_inv0;
  wire [7:0] a0_0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] a0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] b0_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] b0ls1_G4_sq3_G16_inv0_G256_inv0;
  wire [7:0] e0_G16_inv0_G256_inv0;
  wire [7:0] a0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] a0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] b0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] c0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] c0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] d0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] axorb_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] cxord_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] e0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] p0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] q0_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] p0ls1_G4_mul4_G16_inv0_G256_inv0;
  wire [7:0] p0_G16_inv0_G256_inv0;
  wire [7:0] a0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] a0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] b0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] c0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] c0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] d0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] axorb_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] cxord_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] e0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] p0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] q0_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] p0ls1_G4_mul5_G16_inv0_G256_inv0;
  wire [7:0] q0_G16_inv0_G256_inv0;
  wire [7:0] p0ls2_G16_inv0_G256_inv0;
  wire [7:0] e0_G256_inv0;
  wire [7:0] a0_0_G16_mul1_G256_inv0;
  wire [7:0] a0_G16_mul1_G256_inv0;
  wire [7:0] b0_G16_mul1_G256_inv0;
  wire [7:0] c0_0_G16_mul1_G256_inv0;
  wire [7:0] c0_G16_mul1_G256_inv0;
  wire [7:0] d0_G16_mul1_G256_inv0;
  wire [7:0] axorb_0_G16_mul1_G256_inv0;
  wire [7:0] cxord_0_G16_mul1_G256_inv0;
  wire [7:0] a0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] a0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] b0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] c0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] c0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] d0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] axorb_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] cxord_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] e0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] p0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] q0_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] p0ls1_G4_mul0_G16_mul1_G256_inv0;
  wire [7:0] e0_G16_mul1_G256_inv0;
  wire [7:0] a0_0_G4_scl_N0_G16_mul1_G256_inv0;
  wire [7:0] a0_G4_scl_N0_G16_mul1_G256_inv0;
  wire [7:0] b0_G4_scl_N0_G16_mul1_G256_inv0;
  wire [7:0] p0_G4_scl_N0_G16_mul1_G256_inv0;
  wire [7:0] q0_G4_scl_N0_G16_mul1_G256_inv0;
  wire [7:0] p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
  wire [7:0] e01_G16_mul1_G256_inv0;
  wire [7:0] a0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] a0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] b0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] c0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] c0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] d0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] axorb_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] cxord_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] e0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] p0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] q0_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] p0ls1_G4_mul1_G16_mul1_G256_inv0;
  wire [7:0] p0_0_G16_mul1_G256_inv0;
  wire [7:0] p0_G16_mul1_G256_inv0;
  wire [7:0] a0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] a0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] b0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] c0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] c0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] d0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] axorb_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] cxord_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] e0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] p0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] q0_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] p0ls1_G4_mul2_G16_mul1_G256_inv0;
  wire [7:0] q0_0_G16_mul1_G256_inv0;
  wire [7:0] q0_G16_mul1_G256_inv0;
  wire [7:0] p0ls2_G16_mul1_G256_inv0;
  wire [7:0] p0_G256_inv0;
  wire [7:0] a0_0_G16_mul2_G256_inv0;
  wire [7:0] a0_G16_mul2_G256_inv0;
  wire [7:0] b0_G16_mul2_G256_inv0;
  wire [7:0] c0_0_G16_mul2_G256_inv0;
  wire [7:0] c0_G16_mul2_G256_inv0;
  wire [7:0] d0_G16_mul2_G256_inv0;
  wire [7:0] axorb_0_G16_mul2_G256_inv0;
  wire [7:0] cxord_0_G16_mul2_G256_inv0;
  wire [7:0] a0_0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] a0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] b0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] c0_0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] c0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] d0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] axorb_0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] cxord_0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] e0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] p0_0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] p0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] q0_0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] q0_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] p0ls1_G4_mul0_G16_mul2_G256_inv0;
  wire [7:0] e0_G16_mul2_G256_inv0;
  wire [7:0] a0_0_G4_scl_N0_G16_mul2_G256_inv0;
  wire [7:0] a0_G4_scl_N0_G16_mul2_G256_inv0;
  wire [7:0] b0_G4_scl_N0_G16_mul2_G256_inv0;
  wire [7:0] p0_G4_scl_N0_G16_mul2_G256_inv0;
  wire [7:0] q0_G4_scl_N0_G16_mul2_G256_inv0;
  wire [7:0] p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
  wire [7:0] e01_G16_mul2_G256_inv0;
  wire [7:0] a0_0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] a0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] b0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] c0_0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] c0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] d0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] axorb_0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] cxord_0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] e0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] p0_0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] p0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] q0_0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] q0_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] p0ls1_G4_mul1_G16_mul2_G256_inv0;
  wire [7:0] p0_0_G16_mul2_G256_inv0;
  wire [7:0] p0_G16_mul2_G256_inv0;
  wire [7:0] a0_0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] a0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] b0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] c0_0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] c0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] d0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] axorb_0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] cxord_0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] e0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] p0_0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] p0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] q0_0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] q0_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] p0ls1_G4_mul2_G16_mul2_G256_inv0;
  wire [7:0] q0_0_G16_mul2_G256_inv0;
  wire [7:0] q0_G16_mul2_G256_inv0;
  wire [7:0] p0ls2_G16_mul2_G256_inv0;
  wire [7:0] q0_G256_inv0;
  wire [7:0] p0ls4_G256_inv0;
  wire [7:0] t4;
  wire [7:0] y_G256_newbasis1;
  wire [7:0] tempy1_G256_newbasis1;
  wire [7:0] cond1_G256_newbasis1;
  wire [7:0] negCond1_G256_newbasis1;
  wire [7:0] yxorb1_G256_newbasis1;
  wire [7:0] ny1_G256_newbasis1;
  wire [7:0] tempyIntoNegCond1_G256_newbasis1;
  wire [7:0] y1_G256_newbasis1;
  wire [7:0] x1_G256_newbasis1;
  wire [7:0] tempy2_G256_newbasis1;
  wire [7:0] cond2_G256_newbasis1;
  wire [7:0] negCond2_G256_newbasis1;
  wire [7:0] yxorb2_G256_newbasis1;
  wire [7:0] ny2_G256_newbasis1;
  wire [7:0] tempyIntoNegCond2_G256_newbasis1;
  wire [7:0] y2_G256_newbasis1;
  wire [7:0] x2_G256_newbasis1;
  wire [7:0] tempy3_G256_newbasis1;
  wire [7:0] cond3_G256_newbasis1;
  wire [7:0] negCond3_G256_newbasis1;
  wire [7:0] yxorb3_G256_newbasis1;
  wire [7:0] ny3_G256_newbasis1;
  wire [7:0] tempyIntoNegCond3_G256_newbasis1;
  wire [7:0] y3_G256_newbasis1;
  wire [7:0] x3_G256_newbasis1;
  wire [7:0] tempy4_G256_newbasis1;
  wire [7:0] cond4_G256_newbasis1;
  wire [7:0] negCond4_G256_newbasis1;
  wire [7:0] yxorb4_G256_newbasis1;
  wire [7:0] ny4_G256_newbasis1;
  wire [7:0] tempyIntoNegCond4_G256_newbasis1;
  wire [7:0] y4_G256_newbasis1;
  wire [7:0] x4_G256_newbasis1;
  wire [7:0] tempy5_G256_newbasis1;
  wire [7:0] cond5_G256_newbasis1;
  wire [7:0] negCond5_G256_newbasis1;
  wire [7:0] yxorb5_G256_newbasis1;
  wire [7:0] ny5_G256_newbasis1;
  wire [7:0] tempyIntoNegCond5_G256_newbasis1;
  wire [7:0] y5_G256_newbasis1;
  wire [7:0] x5_G256_newbasis1;
  wire [7:0] tempy6_G256_newbasis1;
  wire [7:0] cond6_G256_newbasis1;
  wire [7:0] negCond6_G256_newbasis1;
  wire [7:0] yxorb6_G256_newbasis1;
  wire [7:0] ny6_G256_newbasis1;
  wire [7:0] tempyIntoNegCond6_G256_newbasis1;
  wire [7:0] y6_G256_newbasis1;
  wire [7:0] x6_G256_newbasis1;
  wire [7:0] tempy7_G256_newbasis1;
  wire [7:0] cond7_G256_newbasis1;
  wire [7:0] negCond7_G256_newbasis1;
  wire [7:0] yxorb7_G256_newbasis1;
  wire [7:0] ny7_G256_newbasis1;
  wire [7:0] tempyIntoNegCond7_G256_newbasis1;
  wire [7:0] y7_G256_newbasis1;
  wire [7:0] x7_G256_newbasis1;
  wire [7:0] tempy8_G256_newbasis1;
  wire [7:0] cond8_G256_newbasis1;
  wire [7:0] negCond8_G256_newbasis1;
  wire [7:0] yxorb8_G256_newbasis1;
  wire [7:0] ny8_G256_newbasis1;
  wire [7:0] tempyIntoNegCond8_G256_newbasis1;
  wire [7:0] y8_G256_newbasis1;
  wire [7:0] x8_G256_newbasis1;
  wire [7:0] t6;
  assign dec_99_inp = dec_99;
  assign dec_88_inp = dec_88;
  assign dec_45_inp = dec_45;
  assign dec_158_inp = dec_158;
  assign dec_11_inp = dec_11;
  assign dec_220_inp = dec_220;
  assign dec_36_inp = dec_36;
  assign dec_3_inp = dec_3;
  assign dec_2_inp = dec_2;
  assign dec_12_inp = dec_12;
  assign dec_15_inp = dec_15;
  assign dec_4_inp = dec_4;
  assign dec_240_inp = dec_240;
  assign dec_152_inp = dec_152;
  assign dec_243_inp = dec_243;
  assign dec_242_inp = dec_242;
  assign dec_72_inp = dec_72;
  assign dec_9_inp = dec_9;
  assign dec_129_inp = dec_129;
  assign dec_169_inp = dec_169;
  assign dec_255_inp = dec_255;
  assign dec_1_inp = dec_1;
  assign dec_0_inp = dec_0;
  assign t_inp = t;
  assign y_G256_newbasis0 = dec_0_inp;
  assign tempy1_G256_newbasis0 = y_G256_newbasis0;
  assign cond1_G256_newbasis0 = t_inp & dec_1_inp;
  assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
  assign yxorb1_G256_newbasis0 = y_G256_newbasis0 ^ dec_255_inp;
  assign ny1_G256_newbasis0 = cond1_G256_newbasis0 * yxorb1_G256_newbasis0;
  assign tempyIntoNegCond1_G256_newbasis0 = tempy1_G256_newbasis0 * negCond1_G256_newbasis0;
  assign y1_G256_newbasis0 = ny1_G256_newbasis0 + tempyIntoNegCond1_G256_newbasis0;
  assign x1_G256_newbasis0 = t_inp >> dec_1_inp;
  assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
  assign cond2_G256_newbasis0 = x1_G256_newbasis0 & dec_1_inp;
  assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
  assign yxorb2_G256_newbasis0 = y1_G256_newbasis0 ^ dec_169_inp;
  assign ny2_G256_newbasis0 = cond2_G256_newbasis0 * yxorb2_G256_newbasis0;
  assign tempyIntoNegCond2_G256_newbasis0 = tempy2_G256_newbasis0 * negCond2_G256_newbasis0;
  assign y2_G256_newbasis0 = ny2_G256_newbasis0 + tempyIntoNegCond2_G256_newbasis0;
  assign x2_G256_newbasis0 = x1_G256_newbasis0 >> dec_1_inp;
  assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
  assign cond3_G256_newbasis0 = x2_G256_newbasis0 & dec_1_inp;
  assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
  assign yxorb3_G256_newbasis0 = y2_G256_newbasis0 ^ dec_129_inp;
  assign ny3_G256_newbasis0 = cond3_G256_newbasis0 * yxorb3_G256_newbasis0;
  assign tempyIntoNegCond3_G256_newbasis0 = tempy3_G256_newbasis0 * negCond3_G256_newbasis0;
  assign y3_G256_newbasis0 = ny3_G256_newbasis0 + tempyIntoNegCond3_G256_newbasis0;
  assign x3_G256_newbasis0 = x2_G256_newbasis0 >> dec_1_inp;
  assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
  assign cond4_G256_newbasis0 = x3_G256_newbasis0 & dec_1_inp;
  assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
  assign yxorb4_G256_newbasis0 = y3_G256_newbasis0 ^ dec_9_inp;
  assign ny4_G256_newbasis0 = cond4_G256_newbasis0 * yxorb4_G256_newbasis0;
  assign tempyIntoNegCond4_G256_newbasis0 = tempy4_G256_newbasis0 * negCond4_G256_newbasis0;
  assign y4_G256_newbasis0 = ny4_G256_newbasis0 + tempyIntoNegCond4_G256_newbasis0;
  assign x4_G256_newbasis0 = x3_G256_newbasis0 >> dec_1_inp;
  assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
  assign cond5_G256_newbasis0 = x4_G256_newbasis0 & dec_1_inp;
  assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
  assign yxorb5_G256_newbasis0 = y4_G256_newbasis0 ^ dec_72_inp;
  assign ny5_G256_newbasis0 = cond5_G256_newbasis0 * yxorb5_G256_newbasis0;
  assign tempyIntoNegCond5_G256_newbasis0 = tempy5_G256_newbasis0 * negCond5_G256_newbasis0;
  assign y5_G256_newbasis0 = ny5_G256_newbasis0 + tempyIntoNegCond5_G256_newbasis0;
  assign x5_G256_newbasis0 = x4_G256_newbasis0 >> dec_1_inp;
  assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
  assign cond6_G256_newbasis0 = x5_G256_newbasis0 & dec_1_inp;
  assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
  assign yxorb6_G256_newbasis0 = y5_G256_newbasis0 ^ dec_242_inp;
  assign ny6_G256_newbasis0 = cond6_G256_newbasis0 * yxorb6_G256_newbasis0;
  assign tempyIntoNegCond6_G256_newbasis0 = tempy6_G256_newbasis0 * negCond6_G256_newbasis0;
  assign y6_G256_newbasis0 = ny6_G256_newbasis0 + tempyIntoNegCond6_G256_newbasis0;
  assign x6_G256_newbasis0 = x5_G256_newbasis0 >> dec_1_inp;
  assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
  assign cond7_G256_newbasis0 = x6_G256_newbasis0 & dec_1_inp;
  assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
  assign yxorb7_G256_newbasis0 = y6_G256_newbasis0 ^ dec_243_inp;
  assign ny7_G256_newbasis0 = cond7_G256_newbasis0 * yxorb7_G256_newbasis0;
  assign tempyIntoNegCond7_G256_newbasis0 = tempy7_G256_newbasis0 * negCond7_G256_newbasis0;
  assign y7_G256_newbasis0 = ny7_G256_newbasis0 + tempyIntoNegCond7_G256_newbasis0;
  assign x7_G256_newbasis0 = x6_G256_newbasis0 >> dec_1_inp;
  assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
  assign cond8_G256_newbasis0 = x7_G256_newbasis0 & dec_1_inp;
  assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
  assign yxorb8_G256_newbasis0 = y7_G256_newbasis0 ^ dec_152_inp;
  assign ny8_G256_newbasis0 = cond8_G256_newbasis0 * yxorb8_G256_newbasis0;
  assign tempyIntoNegCond8_G256_newbasis0 = tempy8_G256_newbasis0 * negCond8_G256_newbasis0;
  assign y8_G256_newbasis0 = ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0;
  assign x8_G256_newbasis0 = x7_G256_newbasis0 >> dec_1_inp;
  assign t2 = y8_G256_newbasis0;
  assign a0_0_G256_inv0 = t2 & dec_240_inp;
  assign a0_G256_inv0 = a0_0_G256_inv0 >> dec_4_inp;
  assign b0_G256_inv0 = t2 & dec_15_inp;
  assign a0xorb0_G256_inv0 = a0_G256_inv0 ^ b0_G256_inv0;
  assign a0_0_G16_sq_scl0_G256_inv0 = a0xorb0_G256_inv0 & dec_12_inp;
  assign a0_G16_sq_scl0_G256_inv0 = a0_0_G16_sq_scl0_G256_inv0 >> dec_2_inp;
  assign b0_G16_sq_scl0_G256_inv0 = a0xorb0_G256_inv0 & dec_3_inp;
  assign p0_0_G16_sq_scl0_G256_inv0 = a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0;
  assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = p0_0_G16_sq_scl0_G256_inv0 & dec_2_inp;
  assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp;
  assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = p0_0_G16_sq_scl0_G256_inv0 & dec_1_inp;
  assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = b0_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp;
  assign p0_G16_sq_scl0_G256_inv0 = b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0;
  assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = b0_G16_sq_scl0_G256_inv0 & dec_2_inp;
  assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp;
  assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = b0_G16_sq_scl0_G256_inv0 & dec_1_inp;
  assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = b0_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp;
  assign q0_0_G16_sq_scl0_G256_inv0 = b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0;
  assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = q0_0_G16_sq_scl0_G256_inv0 & dec_2_inp;
  assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp;
  assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = q0_0_G16_sq_scl0_G256_inv0 & dec_1_inp;
  assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp;
  assign q0_G16_sq_scl0_G256_inv0 = p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  assign p0ls2_G16_sq_scl0_G256_inv0 = p0_G16_sq_scl0_G256_inv0 << dec_2_inp;
  assign c0_G256_inv0 = p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0;
  assign a0_0_G16_mul0_G256_inv0 = a0_G256_inv0 & dec_12_inp;
  assign a0_G16_mul0_G256_inv0 = a0_0_G16_mul0_G256_inv0 >> dec_2_inp;
  assign b0_G16_mul0_G256_inv0 = a0_G256_inv0 & dec_3_inp;
  assign c0_0_G16_mul0_G256_inv0 = b0_G256_inv0 & dec_12_inp;
  assign c0_G16_mul0_G256_inv0 = c0_0_G16_mul0_G256_inv0 >> dec_2_inp;
  assign d0_G16_mul0_G256_inv0 = b0_G256_inv0 & dec_3_inp;
  assign axorb_0_G16_mul0_G256_inv0 = a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0;
  assign cxord_0_G16_mul0_G256_inv0 = c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0;
  assign a0_0_G4_mul0_G16_mul0_G256_inv0 = axorb_0_G16_mul0_G256_inv0 & dec_2_inp;
  assign a0_G4_mul0_G16_mul0_G256_inv0 = a0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp;
  assign b0_G4_mul0_G16_mul0_G256_inv0 = axorb_0_G16_mul0_G256_inv0 & dec_1_inp;
  assign c0_0_G4_mul0_G16_mul0_G256_inv0 = cxord_0_G16_mul0_G256_inv0 & dec_2_inp;
  assign c0_G4_mul0_G16_mul0_G256_inv0 = c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul0_G16_mul0_G256_inv0 = cxord_0_G16_mul0_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0;
  assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = c0_G4_mul0_G16_mul0_G256_inv0 ^ d0_G4_mul0_G16_mul0_G256_inv0;
  assign e0_G4_mul0_G16_mul0_G256_inv0 = (dec_243[2])? e0_G4_mul0_G16_mul0_G256_inv0_reg5 & e0_G4_mul0_G16_mul0_G256_inv0_reg6 : ~e0_G4_mul0_G16_mul0_G256_inv0_reg7 & ~e0_G4_mul0_G16_mul0_G256_inv0_reg8;
  assign p0_0_G4_mul0_G16_mul0_G256_inv0 = (dec_12[7])? p0_0_G4_mul0_G16_mul0_G256_inv0_reg1 & p0_0_G4_mul0_G16_mul0_G256_inv0_reg2 : ~p0_0_G4_mul0_G16_mul0_G256_inv0_reg3 & ~p0_0_G4_mul0_G16_mul0_G256_inv0_reg4;
  assign p0_G4_mul0_G16_mul0_G256_inv0 = p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0;
  assign q0_0_G4_mul0_G16_mul0_G256_inv0 = (dec_152[0])? q0_0_G4_mul0_G16_mul0_G256_inv0_reg9 & q0_0_G4_mul0_G16_mul0_G256_inv0_reg10 : ~q0_0_G4_mul0_G16_mul0_G256_inv0_reg11 & ~q0_0_G4_mul0_G16_mul0_G256_inv0_reg12;
  assign q0_G4_mul0_G16_mul0_G256_inv0 = q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0;
  assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = p0_G4_mul0_G16_mul0_G256_inv0 << y_reg122;
  assign e0_G16_mul0_G256_inv0 = p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0;
  assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = e0_G16_mul0_G256_inv0 & y_reg125;
  assign a0_G4_scl_N0_G16_mul0_G256_inv0 = a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> y_reg126;
  assign b0_G4_scl_N0_G16_mul0_G256_inv0 = e0_G16_mul0_G256_inv0 & y_reg123;
  assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
  assign q0_G4_scl_N0_G16_mul0_G256_inv0 = a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0;
  assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = p0_G4_scl_N0_G16_mul0_G256_inv0 << y_reg124;
  assign e01_G16_mul0_G256_inv0 = p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0;
  assign a0_0_G4_mul1_G16_mul0_G256_inv0 = a0_G16_mul0_G256_inv0 & dec_2_inp;
  assign a0_G4_mul1_G16_mul0_G256_inv0 = a0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp;
  assign b0_G4_mul1_G16_mul0_G256_inv0 = a0_G16_mul0_G256_inv0 & dec_1_inp;
  assign c0_0_G4_mul1_G16_mul0_G256_inv0 = c0_G16_mul0_G256_inv0 & dec_2_inp;
  assign c0_G4_mul1_G16_mul0_G256_inv0 = c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul1_G16_mul0_G256_inv0 = c0_G16_mul0_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = e0_G4_mul1_G16_mul0_G256_inv0_reg17 ^ e0_G4_mul1_G16_mul0_G256_inv0_reg18;
  assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = e0_G4_mul1_G16_mul0_G256_inv0_reg19 ^ e0_G4_mul1_G16_mul0_G256_inv0_reg20;
  assign e0_G4_mul1_G16_mul0_G256_inv0 = (dec_9[7])? axorb_0_G4_mul1_G16_mul0_G256_inv0 & cxord_0_G4_mul1_G16_mul0_G256_inv0 : ~e0_G4_mul1_G16_mul0_G256_inv0_reg21 & ~e0_G4_mul1_G16_mul0_G256_inv0_reg22;
  assign p0_0_G4_mul1_G16_mul0_G256_inv0 = (dec_243[5])? p0_0_G4_mul1_G16_mul0_G256_inv0_reg13 & p0_0_G4_mul1_G16_mul0_G256_inv0_reg14 : ~p0_0_G4_mul1_G16_mul0_G256_inv0_reg15 & ~p0_0_G4_mul1_G16_mul0_G256_inv0_reg16;
  assign p0_G4_mul1_G16_mul0_G256_inv0 = p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0;
  assign q0_0_G4_mul1_G16_mul0_G256_inv0 = (dec_243[6])? q0_0_G4_mul1_G16_mul0_G256_inv0_reg23 & q0_0_G4_mul1_G16_mul0_G256_inv0_reg24 : ~q0_0_G4_mul1_G16_mul0_G256_inv0_reg25 & ~q0_0_G4_mul1_G16_mul0_G256_inv0_reg26;
  assign q0_G4_mul1_G16_mul0_G256_inv0 = q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0;
  assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = p0_G4_mul1_G16_mul0_G256_inv0 << y_reg121;
  assign p0_0_G16_mul0_G256_inv0 = p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0;
  assign p0_G16_mul0_G256_inv0 = p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0;
  assign a0_0_G4_mul2_G16_mul0_G256_inv0 = b0_G16_mul0_G256_inv0 & dec_2_inp;
  assign a0_G4_mul2_G16_mul0_G256_inv0 = a0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp;
  assign b0_G4_mul2_G16_mul0_G256_inv0 = b0_G16_mul0_G256_inv0 & dec_1_inp;
  assign c0_0_G4_mul2_G16_mul0_G256_inv0 = d0_G16_mul0_G256_inv0 & dec_2_inp;
  assign c0_G4_mul2_G16_mul0_G256_inv0 = c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul2_G16_mul0_G256_inv0 = d0_G16_mul0_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = e0_G4_mul2_G16_mul0_G256_inv0_reg31 ^ e0_G4_mul2_G16_mul0_G256_inv0_reg32;
  assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = e0_G4_mul2_G16_mul0_G256_inv0_reg33 ^ e0_G4_mul2_G16_mul0_G256_inv0_reg34;
  assign e0_G4_mul2_G16_mul0_G256_inv0 = (dec_0[5])? axorb_0_G4_mul2_G16_mul0_G256_inv0 & cxord_0_G4_mul2_G16_mul0_G256_inv0 : ~e0_G4_mul2_G16_mul0_G256_inv0_reg35 & ~e0_G4_mul2_G16_mul0_G256_inv0_reg36;
  assign p0_0_G4_mul2_G16_mul0_G256_inv0 = (dec_12[0])? p0_0_G4_mul2_G16_mul0_G256_inv0_reg27 & p0_0_G4_mul2_G16_mul0_G256_inv0_reg28 : p0_0_G4_mul2_G16_mul0_G256_inv0_reg29 & p0_0_G4_mul2_G16_mul0_G256_inv0_reg30;
  assign p0_G4_mul2_G16_mul0_G256_inv0 = p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0;
  assign q0_0_G4_mul2_G16_mul0_G256_inv0 = (dec_169[1])? q0_0_G4_mul2_G16_mul0_G256_inv0_reg37 & q0_0_G4_mul2_G16_mul0_G256_inv0_reg38 : ~q0_0_G4_mul2_G16_mul0_G256_inv0_reg39 & ~q0_0_G4_mul2_G16_mul0_G256_inv0_reg40;
  assign q0_G4_mul2_G16_mul0_G256_inv0 = q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0;
  assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = p0_G4_mul2_G16_mul0_G256_inv0 << y_reg128;
  assign q0_0_G16_mul0_G256_inv0 = p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0;
  assign q0_G16_mul0_G256_inv0 = q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0;
  assign p0ls2_G16_mul0_G256_inv0 = p0_G16_mul0_G256_inv0 << y_reg127;
  assign d0_G256_inv0 = p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0;
  assign c0xord0_G256_inv0 = y_reg129 ^ d0_G256_inv0;
  assign a0_0_G16_inv0_G256_inv0 = c0xord0_G256_inv0 & y_reg130;
  assign a0_G16_inv0_G256_inv0 = a0_0_G16_inv0_G256_inv0 >> y_reg131;
  assign b0_G16_inv0_G256_inv0 = c0xord0_G256_inv0 & y_reg132;
  assign a0xorb0_G16_inv0_G256_inv0 = a0_G16_inv0_G256_inv0 ^ b0_G16_inv0_G256_inv0;
  assign a0_0_G4_sq2_G16_inv0_G256_inv0 = a0xorb0_G16_inv0_G256_inv0 & y_reg135;
  assign a0_G4_sq2_G16_inv0_G256_inv0 = a0_0_G4_sq2_G16_inv0_G256_inv0 >> y_reg136;
  assign b0_G4_sq2_G16_inv0_G256_inv0 = a0xorb0_G16_inv0_G256_inv0 & y_reg133;
  assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = b0_G4_sq2_G16_inv0_G256_inv0 << y_reg134;
  assign c0_0_G16_inv0_G256_inv0 = b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0;
  assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = c0_0_G16_inv0_G256_inv0 & y_reg139;
  assign a0_G4_scl_N1_G16_inv0_G256_inv0 = a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> y_reg140;
  assign b0_G4_scl_N1_G16_inv0_G256_inv0 = c0_0_G16_inv0_G256_inv0 & y_reg137;
  assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
  assign q0_G4_scl_N1_G16_inv0_G256_inv0 = a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0;
  assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = p0_G4_scl_N1_G16_inv0_G256_inv0 << y_reg138;
  assign c0_G16_inv0_G256_inv0 = p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0;
  assign a0_0_G4_mul3_G16_inv0_G256_inv0 = a0_G16_inv0_G256_inv0 & y_reg150;
  assign a0_G4_mul3_G16_inv0_G256_inv0 = a0_0_G4_mul3_G16_inv0_G256_inv0 >> y_reg151;
  assign b0_G4_mul3_G16_inv0_G256_inv0 = a0_G16_inv0_G256_inv0 & y_reg169;
  assign c0_0_G4_mul3_G16_inv0_G256_inv0 = b0_G16_inv0_G256_inv0 & y_reg152;
  assign c0_G4_mul3_G16_inv0_G256_inv0 = c0_0_G4_mul3_G16_inv0_G256_inv0 >> y_reg153;
  assign d0_G4_mul3_G16_inv0_G256_inv0 = b0_G16_inv0_G256_inv0 & y_reg170;
  assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = e0_G4_mul3_G16_inv0_G256_inv0_reg45 ^ e0_G4_mul3_G16_inv0_G256_inv0_reg46;
  assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = e0_G4_mul3_G16_inv0_G256_inv0_reg47 ^ e0_G4_mul3_G16_inv0_G256_inv0_reg48;
  assign e0_G4_mul3_G16_inv0_G256_inv0 = (r[13])? axorb_0_G4_mul3_G16_inv0_G256_inv0 & cxord_0_G4_mul3_G16_inv0_G256_inv0 : e0_G4_mul3_G16_inv0_G256_inv0_reg49 & e0_G4_mul3_G16_inv0_G256_inv0_reg50;
  assign p0_0_G4_mul3_G16_inv0_G256_inv0 = (dec_36[5])? p0_0_G4_mul3_G16_inv0_G256_inv0_reg41 & p0_0_G4_mul3_G16_inv0_G256_inv0_reg42 : p0_0_G4_mul3_G16_inv0_G256_inv0_reg43 & p0_0_G4_mul3_G16_inv0_G256_inv0_reg44;
  assign p0_G4_mul3_G16_inv0_G256_inv0 = p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0;
  assign q0_0_G4_mul3_G16_inv0_G256_inv0 = (dec_242[4])? q0_0_G4_mul3_G16_inv0_G256_inv0_reg51 & q0_0_G4_mul3_G16_inv0_G256_inv0_reg52 : ~q0_0_G4_mul3_G16_inv0_G256_inv0_reg53 & ~q0_0_G4_mul3_G16_inv0_G256_inv0_reg54;
  assign q0_G4_mul3_G16_inv0_G256_inv0 = q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0;
  assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = p0_G4_mul3_G16_inv0_G256_inv0 << y_reg172;
  assign d0_G16_inv0_G256_inv0 = p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0;
  assign c0xord0_G16_inv0_G256_inv0 = y_reg181 ^ d0_G16_inv0_G256_inv0;
  assign a0_0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg204;
  assign a0_G4_sq3_G16_inv0_G256_inv0 = a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg206;
  assign b0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg200;
  assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = b0_G4_sq3_G16_inv0_G256_inv0 << y_reg202;
  assign e0_G16_inv0_G256_inv0 = b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0;
  assign a0_0_G4_mul4_G16_inv0_G256_inv0 = e0_G16_inv0_G256_inv0 & y_reg208;
  assign a0_G4_mul4_G16_inv0_G256_inv0 = a0_0_G4_mul4_G16_inv0_G256_inv0 >> y_reg210;
  assign b0_G4_mul4_G16_inv0_G256_inv0 = e0_G16_inv0_G256_inv0 & y_reg241;
  assign c0_0_G4_mul4_G16_inv0_G256_inv0 = b0_G16_inv0_G256_inv0 & y_reg211;
  assign c0_G4_mul4_G16_inv0_G256_inv0 = c0_0_G4_mul4_G16_inv0_G256_inv0 >> y_reg212;
  assign d0_G4_mul4_G16_inv0_G256_inv0 = b0_G16_inv0_G256_inv0 & y_reg242;
  assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0;
  assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = c0_G4_mul4_G16_inv0_G256_inv0 ^ d0_G4_mul4_G16_inv0_G256_inv0;
  assign e0_G4_mul4_G16_inv0_G256_inv0 = (dec_255[0])? e0_G4_mul4_G16_inv0_G256_inv0_reg59 & y_reg243 : ~e0_G4_mul4_G16_inv0_G256_inv0_reg61 & y_reg239;
  assign p0_0_G4_mul4_G16_inv0_G256_inv0 = (t[4])? p0_0_G4_mul4_G16_inv0_G256_inv0_reg55 & y_reg213 : ~p0_0_G4_mul4_G16_inv0_G256_inv0_reg57 & y_reg198;
  assign p0_G4_mul4_G16_inv0_G256_inv0 = p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0;
  assign q0_0_G4_mul4_G16_inv0_G256_inv0 = (dec_45[1])? q0_0_G4_mul4_G16_inv0_G256_inv0_reg63 & y_reg264 : ~q0_0_G4_mul4_G16_inv0_G256_inv0_reg65 & y_reg263;
  assign q0_G4_mul4_G16_inv0_G256_inv0 = q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0;
  assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = p0_G4_mul4_G16_inv0_G256_inv0 << y_reg246;
  assign p0_G16_inv0_G256_inv0 = p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0;
  assign a0_0_G4_mul5_G16_inv0_G256_inv0 = e0_G16_inv0_G256_inv0 & y_reg287;
  assign a0_G4_mul5_G16_inv0_G256_inv0 = a0_0_G4_mul5_G16_inv0_G256_inv0 >> y_reg289;
  assign b0_G4_mul5_G16_inv0_G256_inv0 = e0_G16_inv0_G256_inv0 & y_reg321;
  assign c0_0_G4_mul5_G16_inv0_G256_inv0 = a0_G16_inv0_G256_inv0 & y_reg290;
  assign c0_G4_mul5_G16_inv0_G256_inv0 = c0_0_G4_mul5_G16_inv0_G256_inv0 >> y_reg291;
  assign d0_G4_mul5_G16_inv0_G256_inv0 = a0_G16_inv0_G256_inv0 & y_reg322;
  assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = e0_G4_mul5_G16_inv0_G256_inv0_reg71 ^ e0_G4_mul5_G16_inv0_G256_inv0_reg72;
  assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = e0_G4_mul5_G16_inv0_G256_inv0_reg73 ^ e0_G4_mul5_G16_inv0_G256_inv0_reg74;
  assign e0_G4_mul5_G16_inv0_G256_inv0 = (dec_3[1])? axorb_0_G4_mul5_G16_inv0_G256_inv0 & y_reg323 : ~e0_G4_mul5_G16_inv0_G256_inv0_reg75 & y_reg319;
  assign p0_0_G4_mul5_G16_inv0_G256_inv0 = (dec_99[0])? p0_0_G4_mul5_G16_inv0_G256_inv0_reg67 & y_reg292 : ~p0_0_G4_mul5_G16_inv0_G256_inv0_reg69 & y_reg285;
  assign p0_G4_mul5_G16_inv0_G256_inv0 = p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0;
  assign q0_0_G4_mul5_G16_inv0_G256_inv0 = (dec_9[1])? q0_0_G4_mul5_G16_inv0_G256_inv0_reg77 & y_reg344 : ~q0_0_G4_mul5_G16_inv0_G256_inv0_reg79 & y_reg343;
  assign q0_G4_mul5_G16_inv0_G256_inv0 = q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0;
  assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = p0_G4_mul5_G16_inv0_G256_inv0 << y_reg326;
  assign q0_G16_inv0_G256_inv0 = p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0;
  assign p0ls2_G16_inv0_G256_inv0 = p0_G16_inv0_G256_inv0 << y_reg267;
  assign e0_G256_inv0 = p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0;
  assign a0_0_G16_mul1_G256_inv0 = e0_G256_inv0 & y_reg362;
  assign a0_G16_mul1_G256_inv0 = a0_0_G16_mul1_G256_inv0 >> y_reg365;
  assign b0_G16_mul1_G256_inv0 = e0_G256_inv0 & y_reg447;
  assign c0_0_G16_mul1_G256_inv0 = b0_G256_inv0 & dec_12_inp;
  assign c0_G16_mul1_G256_inv0 = c0_0_G16_mul1_G256_inv0 >> dec_2_inp;
  assign d0_G16_mul1_G256_inv0 = b0_G256_inv0 & dec_3_inp;
  assign axorb_0_G16_mul1_G256_inv0 = a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0;
  assign cxord_0_G16_mul1_G256_inv0 = c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0;
  assign a0_0_G4_mul0_G16_mul1_G256_inv0 = axorb_0_G16_mul1_G256_inv0 & y_reg450;
  assign a0_G4_mul0_G16_mul1_G256_inv0 = a0_0_G4_mul0_G16_mul1_G256_inv0 >> y_reg453;
  assign b0_G4_mul0_G16_mul1_G256_inv0 = axorb_0_G16_mul1_G256_inv0 & y_reg486;
  assign c0_0_G4_mul0_G16_mul1_G256_inv0 = cxord_0_G16_mul1_G256_inv0 & dec_2_inp;
  assign c0_G4_mul0_G16_mul1_G256_inv0 = c0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul0_G16_mul1_G256_inv0 = cxord_0_G16_mul1_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = e0_G4_mul0_G16_mul1_G256_inv0_reg85 ^ e0_G4_mul0_G16_mul1_G256_inv0_reg86;
  assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = e0_G4_mul0_G16_mul1_G256_inv0_reg87 ^ e0_G4_mul0_G16_mul1_G256_inv0_reg88;
  assign e0_G4_mul0_G16_mul1_G256_inv0 = (dec_36[7])? axorb_0_G4_mul0_G16_mul1_G256_inv0 & y_reg489 : ~e0_G4_mul0_G16_mul1_G256_inv0_reg89 & y_reg483;
  assign p0_0_G4_mul0_G16_mul1_G256_inv0 = (dec_11[2])? p0_0_G4_mul0_G16_mul1_G256_inv0_reg81 & y_reg456 : ~p0_0_G4_mul0_G16_mul1_G256_inv0_reg83 & y_reg444;
  assign p0_G4_mul0_G16_mul1_G256_inv0 = p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0;
  assign q0_0_G4_mul0_G16_mul1_G256_inv0 = (dec_12[3])? q0_0_G4_mul0_G16_mul1_G256_inv0_reg91 & y_reg514 : q0_0_G4_mul0_G16_mul1_G256_inv0_reg93 & y_reg511;
  assign q0_G4_mul0_G16_mul1_G256_inv0 = q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0;
  assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = p0_G4_mul0_G16_mul1_G256_inv0 << y_reg493;
  assign e0_G16_mul1_G256_inv0 = p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0;
  assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = e0_G16_mul1_G256_inv0 & y_reg526;
  assign a0_G4_scl_N0_G16_mul1_G256_inv0 = a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> y_reg530;
  assign b0_G4_scl_N0_G16_mul1_G256_inv0 = e0_G16_mul1_G256_inv0 & y_reg518;
  assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
  assign q0_G4_scl_N0_G16_mul1_G256_inv0 = a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0;
  assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = p0_G4_scl_N0_G16_mul1_G256_inv0 << y_reg522;
  assign e01_G16_mul1_G256_inv0 = p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0;
  assign a0_0_G4_mul1_G16_mul1_G256_inv0 = a0_G16_mul1_G256_inv0 & y_reg368;
  assign a0_G4_mul1_G16_mul1_G256_inv0 = a0_0_G4_mul1_G16_mul1_G256_inv0 >> y_reg371;
  assign b0_G4_mul1_G16_mul1_G256_inv0 = a0_G16_mul1_G256_inv0 & y_reg401;
  assign c0_0_G4_mul1_G16_mul1_G256_inv0 = c0_G16_mul1_G256_inv0 & dec_2_inp;
  assign c0_G4_mul1_G16_mul1_G256_inv0 = c0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul1_G16_mul1_G256_inv0 = c0_G16_mul1_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = e0_G4_mul1_G16_mul1_G256_inv0_reg99 ^ e0_G4_mul1_G16_mul1_G256_inv0_reg100;
  assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = e0_G4_mul1_G16_mul1_G256_inv0_reg101 ^ e0_G4_mul1_G16_mul1_G256_inv0_reg102;
  assign e0_G4_mul1_G16_mul1_G256_inv0 = (dec_88[0])? axorb_0_G4_mul1_G16_mul1_G256_inv0 & y_reg404 : ~e0_G4_mul1_G16_mul1_G256_inv0_reg103 & y_reg398;
  assign p0_0_G4_mul1_G16_mul1_G256_inv0 = (dec_1[1])? p0_0_G4_mul1_G16_mul1_G256_inv0_reg95 & y_reg374 : ~p0_0_G4_mul1_G16_mul1_G256_inv0_reg97 & y_reg359;
  assign p0_G4_mul1_G16_mul1_G256_inv0 = p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0;
  assign q0_0_G4_mul1_G16_mul1_G256_inv0 = (dec_3[1])? q0_0_G4_mul1_G16_mul1_G256_inv0_reg105 & y_reg426 : ~q0_0_G4_mul1_G16_mul1_G256_inv0_reg107 & y_reg423;
  assign q0_G4_mul1_G16_mul1_G256_inv0 = q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0;
  assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = p0_G4_mul1_G16_mul1_G256_inv0 << y_reg408;
  assign p0_0_G16_mul1_G256_inv0 = p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0;
  assign p0_G16_mul1_G256_inv0 = p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0;
  assign a0_0_G4_mul2_G16_mul1_G256_inv0 = b0_G16_mul1_G256_inv0 & y_reg552;
  assign a0_G4_mul2_G16_mul1_G256_inv0 = a0_0_G4_mul2_G16_mul1_G256_inv0 >> y_reg555;
  assign b0_G4_mul2_G16_mul1_G256_inv0 = b0_G16_mul1_G256_inv0 & y_reg582;
  assign c0_0_G4_mul2_G16_mul1_G256_inv0 = d0_G16_mul1_G256_inv0 & dec_2_inp;
  assign c0_G4_mul2_G16_mul1_G256_inv0 = c0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul2_G16_mul1_G256_inv0 = d0_G16_mul1_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0;
  assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = c0_G4_mul2_G16_mul1_G256_inv0 ^ d0_G4_mul2_G16_mul1_G256_inv0;
  assign e0_G4_mul2_G16_mul1_G256_inv0 = (dec_11[2])? e0_G4_mul2_G16_mul1_G256_inv0_reg113 & y_reg585 : ~e0_G4_mul2_G16_mul1_G256_inv0_reg115 & y_reg579;
  assign p0_0_G4_mul2_G16_mul1_G256_inv0 = (r[19])? p0_0_G4_mul2_G16_mul1_G256_inv0_reg109 & y_reg558 : ~p0_0_G4_mul2_G16_mul1_G256_inv0_reg111 & y_reg549;
  assign p0_G4_mul2_G16_mul1_G256_inv0 = p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0;
  assign q0_0_G4_mul2_G16_mul1_G256_inv0 = (dec_72[7])? q0_0_G4_mul2_G16_mul1_G256_inv0_reg117 & y_reg607 : ~q0_0_G4_mul2_G16_mul1_G256_inv0_reg119 & y_reg604;
  assign q0_G4_mul2_G16_mul1_G256_inv0 = q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0;
  assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = p0_G4_mul2_G16_mul1_G256_inv0 << y_reg589;
  assign q0_0_G16_mul1_G256_inv0 = p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0;
  assign q0_G16_mul1_G256_inv0 = q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0;
  assign p0ls2_G16_mul1_G256_inv0 = p0_G16_mul1_G256_inv0 << y_reg534;
  assign p0_G256_inv0 = p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0;
  assign a0_0_G16_mul2_G256_inv0 = e0_G256_inv0 & y_reg614;
  assign a0_G16_mul2_G256_inv0 = a0_0_G16_mul2_G256_inv0 >> y_reg617;
  assign b0_G16_mul2_G256_inv0 = e0_G256_inv0 & y_reg641;
  assign c0_0_G16_mul2_G256_inv0 = a0_G256_inv0 & dec_12_inp;
  assign c0_G16_mul2_G256_inv0 = c0_0_G16_mul2_G256_inv0 >> dec_2_inp;
  assign d0_G16_mul2_G256_inv0 = a0_G256_inv0 & dec_3_inp;
  assign axorb_0_G16_mul2_G256_inv0 = a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0;
  assign cxord_0_G16_mul2_G256_inv0 = c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0;
  assign a0_0_G4_mul0_G16_mul2_G256_inv0 = axorb_0_G16_mul2_G256_inv0 & y_reg644;
  assign a0_G4_mul0_G16_mul2_G256_inv0 = a0_0_G4_mul0_G16_mul2_G256_inv0 >> y_reg647;
  assign b0_G4_mul0_G16_mul2_G256_inv0 = axorb_0_G16_mul2_G256_inv0 & y_reg653;
  assign c0_0_G4_mul0_G16_mul2_G256_inv0 = cxord_0_G16_mul2_G256_inv0 & dec_2_inp;
  assign c0_G4_mul0_G16_mul2_G256_inv0 = c0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul0_G16_mul2_G256_inv0 = cxord_0_G16_mul2_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0;
  assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = c0_G4_mul0_G16_mul2_G256_inv0 ^ d0_G4_mul0_G16_mul2_G256_inv0;
  assign e0_G4_mul0_G16_mul2_G256_inv0 = axorb_0_G4_mul0_G16_mul2_G256_inv0 & y_reg656;
  assign p0_0_G4_mul0_G16_mul2_G256_inv0 = a0_G4_mul0_G16_mul2_G256_inv0 & y_reg650;
  assign p0_G4_mul0_G16_mul2_G256_inv0 = p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0;
  assign q0_0_G4_mul0_G16_mul2_G256_inv0 = b0_G4_mul0_G16_mul2_G256_inv0 & y_reg662;
  assign q0_G4_mul0_G16_mul2_G256_inv0 = q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0;
  assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = p0_G4_mul0_G16_mul2_G256_inv0 << y_reg659;
  assign e0_G16_mul2_G256_inv0 = p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0;
  assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = e0_G16_mul2_G256_inv0 & y_reg671;
  assign a0_G4_scl_N0_G16_mul2_G256_inv0 = a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> y_reg674;
  assign b0_G4_scl_N0_G16_mul2_G256_inv0 = e0_G16_mul2_G256_inv0 & y_reg665;
  assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
  assign q0_G4_scl_N0_G16_mul2_G256_inv0 = a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0;
  assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = p0_G4_scl_N0_G16_mul2_G256_inv0 << y_reg668;
  assign e01_G16_mul2_G256_inv0 = p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0;
  assign a0_0_G4_mul1_G16_mul2_G256_inv0 = a0_G16_mul2_G256_inv0 & y_reg620;
  assign a0_G4_mul1_G16_mul2_G256_inv0 = a0_0_G4_mul1_G16_mul2_G256_inv0 >> y_reg623;
  assign b0_G4_mul1_G16_mul2_G256_inv0 = a0_G16_mul2_G256_inv0 & y_reg629;
  assign c0_0_G4_mul1_G16_mul2_G256_inv0 = c0_G16_mul2_G256_inv0 & dec_2_inp;
  assign c0_G4_mul1_G16_mul2_G256_inv0 = c0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul1_G16_mul2_G256_inv0 = c0_G16_mul2_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0;
  assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = c0_G4_mul1_G16_mul2_G256_inv0 ^ d0_G4_mul1_G16_mul2_G256_inv0;
  assign e0_G4_mul1_G16_mul2_G256_inv0 = axorb_0_G4_mul1_G16_mul2_G256_inv0 & y_reg632;
  assign p0_0_G4_mul1_G16_mul2_G256_inv0 = a0_G4_mul1_G16_mul2_G256_inv0 & y_reg626;
  assign p0_G4_mul1_G16_mul2_G256_inv0 = p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0;
  assign q0_0_G4_mul1_G16_mul2_G256_inv0 = b0_G4_mul1_G16_mul2_G256_inv0 & y_reg638;
  assign q0_G4_mul1_G16_mul2_G256_inv0 = q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0;
  assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = p0_G4_mul1_G16_mul2_G256_inv0 << y_reg635;
  assign p0_0_G16_mul2_G256_inv0 = p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0;
  assign p0_G16_mul2_G256_inv0 = p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0;
  assign a0_0_G4_mul2_G16_mul2_G256_inv0 = b0_G16_mul2_G256_inv0 & y_reg680;
  assign a0_G4_mul2_G16_mul2_G256_inv0 = a0_0_G4_mul2_G16_mul2_G256_inv0 >> y_reg683;
  assign b0_G4_mul2_G16_mul2_G256_inv0 = b0_G16_mul2_G256_inv0 & y_reg689;
  assign c0_0_G4_mul2_G16_mul2_G256_inv0 = d0_G16_mul2_G256_inv0 & dec_2_inp;
  assign c0_G4_mul2_G16_mul2_G256_inv0 = c0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp;
  assign d0_G4_mul2_G16_mul2_G256_inv0 = d0_G16_mul2_G256_inv0 & dec_1_inp;
  assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0;
  assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = c0_G4_mul2_G16_mul2_G256_inv0 ^ d0_G4_mul2_G16_mul2_G256_inv0;
  assign e0_G4_mul2_G16_mul2_G256_inv0 = axorb_0_G4_mul2_G16_mul2_G256_inv0 & y_reg692;
  assign p0_0_G4_mul2_G16_mul2_G256_inv0 = a0_G4_mul2_G16_mul2_G256_inv0 & y_reg686;
  assign p0_G4_mul2_G16_mul2_G256_inv0 = p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0;
  assign q0_0_G4_mul2_G16_mul2_G256_inv0 = b0_G4_mul2_G16_mul2_G256_inv0 & y_reg698;
  assign q0_G4_mul2_G16_mul2_G256_inv0 = q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0;
  assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = p0_G4_mul2_G16_mul2_G256_inv0 << y_reg695;
  assign q0_0_G16_mul2_G256_inv0 = p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0;
  assign q0_G16_mul2_G256_inv0 = q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0;
  assign p0ls2_G16_mul2_G256_inv0 = p0_G16_mul2_G256_inv0 << y_reg677;
  assign q0_G256_inv0 = p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0;
  assign p0ls4_G256_inv0 = p0_G256_inv0 << y_reg611;
  assign t4 = p0ls4_G256_inv0 | y_reg699;
  assign y_G256_newbasis1 = dec_0_inp;
  assign tempy1_G256_newbasis1 = y_G256_newbasis1;
  assign cond1_G256_newbasis1 = t4 & y_reg759;
  assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
  assign yxorb1_G256_newbasis1 = y_G256_newbasis1 ^ dec_36_inp;
  assign ny1_G256_newbasis1 = cond1_G256_newbasis1 * y_reg763;
  assign tempyIntoNegCond1_G256_newbasis1 = y_reg767 * negCond1_G256_newbasis1;
  assign y1_G256_newbasis1 = ny1_G256_newbasis1 + tempyIntoNegCond1_G256_newbasis1;
  assign x1_G256_newbasis1 = t4 >> y_reg703;
  assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
  assign cond2_G256_newbasis1 = x1_G256_newbasis1 & y_reg755;
  assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
  assign yxorb2_G256_newbasis1 = y1_G256_newbasis1 ^ y_reg771;
  assign ny2_G256_newbasis1 = cond2_G256_newbasis1 * yxorb2_G256_newbasis1;
  assign tempyIntoNegCond2_G256_newbasis1 = tempy2_G256_newbasis1 * negCond2_G256_newbasis1;
  assign y2_G256_newbasis1 = ny2_G256_newbasis1 + tempyIntoNegCond2_G256_newbasis1;
  assign x2_G256_newbasis1 = x1_G256_newbasis1 >> y_reg707;
  assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
  assign cond3_G256_newbasis1 = x2_G256_newbasis1 & y_reg751;
  assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
  assign yxorb3_G256_newbasis1 = y2_G256_newbasis1 ^ y_reg775;
  assign ny3_G256_newbasis1 = cond3_G256_newbasis1 * yxorb3_G256_newbasis1;
  assign tempyIntoNegCond3_G256_newbasis1 = tempy3_G256_newbasis1 * negCond3_G256_newbasis1;
  assign y3_G256_newbasis1 = ny3_G256_newbasis1 + tempyIntoNegCond3_G256_newbasis1;
  assign x3_G256_newbasis1 = x2_G256_newbasis1 >> y_reg711;
  assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
  assign cond4_G256_newbasis1 = x3_G256_newbasis1 & y_reg747;
  assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
  assign yxorb4_G256_newbasis1 = y3_G256_newbasis1 ^ y_reg779;
  assign ny4_G256_newbasis1 = cond4_G256_newbasis1 * yxorb4_G256_newbasis1;
  assign tempyIntoNegCond4_G256_newbasis1 = tempy4_G256_newbasis1 * negCond4_G256_newbasis1;
  assign y4_G256_newbasis1 = ny4_G256_newbasis1 + tempyIntoNegCond4_G256_newbasis1;
  assign x4_G256_newbasis1 = x3_G256_newbasis1 >> y_reg715;
  assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
  assign cond5_G256_newbasis1 = x4_G256_newbasis1 & y_reg743;
  assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
  assign yxorb5_G256_newbasis1 = y4_G256_newbasis1 ^ y_reg783;
  assign ny5_G256_newbasis1 = cond5_G256_newbasis1 * yxorb5_G256_newbasis1;
  assign tempyIntoNegCond5_G256_newbasis1 = tempy5_G256_newbasis1 * negCond5_G256_newbasis1;
  assign y5_G256_newbasis1 = ny5_G256_newbasis1 + tempyIntoNegCond5_G256_newbasis1;
  assign x5_G256_newbasis1 = x4_G256_newbasis1 >> y_reg719;
  assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
  assign cond6_G256_newbasis1 = x5_G256_newbasis1 & y_reg739;
  assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
  assign yxorb6_G256_newbasis1 = y5_G256_newbasis1 ^ y_reg787;
  assign ny6_G256_newbasis1 = cond6_G256_newbasis1 * yxorb6_G256_newbasis1;
  assign tempyIntoNegCond6_G256_newbasis1 = tempy6_G256_newbasis1 * negCond6_G256_newbasis1;
  assign y6_G256_newbasis1 = ny6_G256_newbasis1 + tempyIntoNegCond6_G256_newbasis1;
  assign x6_G256_newbasis1 = x5_G256_newbasis1 >> y_reg723;
  assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
  assign cond7_G256_newbasis1 = x6_G256_newbasis1 & y_reg735;
  assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
  assign yxorb7_G256_newbasis1 = y6_G256_newbasis1 ^ y_reg791;
  assign ny7_G256_newbasis1 = cond7_G256_newbasis1 * yxorb7_G256_newbasis1;
  assign tempyIntoNegCond7_G256_newbasis1 = tempy7_G256_newbasis1 * negCond7_G256_newbasis1;
  assign y7_G256_newbasis1 = ny7_G256_newbasis1 + tempyIntoNegCond7_G256_newbasis1;
  assign x7_G256_newbasis1 = x6_G256_newbasis1 >> y_reg727;
  assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
  assign cond8_G256_newbasis1 = x7_G256_newbasis1 & y_reg731;
  assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
  assign yxorb8_G256_newbasis1 = y7_G256_newbasis1 ^ y_reg795;
  assign ny8_G256_newbasis1 = cond8_G256_newbasis1 * yxorb8_G256_newbasis1;
  assign tempyIntoNegCond8_G256_newbasis1 = tempy8_G256_newbasis1 * negCond8_G256_newbasis1;
  assign y8_G256_newbasis1 = ny8_G256_newbasis1 + tempyIntoNegCond8_G256_newbasis1;
  assign x8_G256_newbasis1 = x7_G256_newbasis1 >> dec_1_inp;
  assign t6 = y8_G256_newbasis1;

  always @(posedge clk) begin
    y <= t6 ^ y_reg799;
  end

  assign t5_a0_0_G16_mul0_G256_inv0 = ~(~a0_G256_inv0 | ~dec_12_inp);
  assign t6_dec_2_inp = dec_2;
  assign t4_a0_G16_mul0_G256_inv0 = t5_a0_0_G16_mul0_G256_inv0 >> t6_dec_2_inp;
  assign t8_a0_G256_inv0 = a0_0_G256_inv0 >> dec_4_inp;
  assign t9_dec_3_inp = ~(~dec_3);
  assign t7_b0_G16_mul0_G256_inv0 = t8_a0_G256_inv0 & t9_dec_3_inp;
  assign t3_axorb_0_G16_mul0_G256_inv0 = ~(~t4_a0_G16_mul0_G256_inv0 ^ t7_b0_G16_mul0_G256_inv0);
  assign t10_dec_2_inp = dec_2;
  assign t2_a0_0_G4_mul0_G16_mul0_G256_inv0 = ~(~t3_axorb_0_G16_mul0_G256_inv0 | ~t10_dec_2_inp);
  assign t11_dec_1_inp = dec_1;
  assign t1_a0_G4_mul0_G16_mul0_G256_inv0 = ~(t2_a0_0_G4_mul0_G16_mul0_G256_inv0 >> t11_dec_1_inp);
  assign t16_c0_0_G16_mul0_G256_inv0 = b0_G256_inv0 & dec_12_inp;
  assign t17_dec_2_inp = dec_2;
  assign t15_c0_G16_mul0_G256_inv0 = ~(~(t16_c0_0_G16_mul0_G256_inv0 >> t17_dec_2_inp));
  assign t19_b0_G256_inv0 = ~(~t2 | ~dec_15_inp);
  assign t20_dec_3_inp = ~(~dec_3);
  assign t18_d0_G16_mul0_G256_inv0 = ~(~t19_b0_G256_inv0 | ~t20_dec_3_inp);
  assign t14_cxord_0_G16_mul0_G256_inv0 = t15_c0_G16_mul0_G256_inv0 ^ t18_d0_G16_mul0_G256_inv0;
  assign t21_dec_2_inp = ~(~dec_2);
  assign t13_c0_0_G4_mul0_G16_mul0_G256_inv0 = t14_cxord_0_G16_mul0_G256_inv0 & t21_dec_2_inp;
  assign t22_dec_1_inp = dec_1;
  assign t12_c0_G4_mul0_G16_mul0_G256_inv0 = ~(t13_c0_0_G4_mul0_G16_mul0_G256_inv0 >> t22_dec_1_inp);
  wire clk1;
  assign clk1 = dec_12[7] & clk;

  always @(posedge clk1) begin
    p0_0_G4_mul0_G16_mul0_G256_inv0_reg1 <= a0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk2;
  assign clk2 = dec_12[7] & clk;

  always @(posedge clk2) begin
    p0_0_G4_mul0_G16_mul0_G256_inv0_reg2 <= c0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk3;
  assign clk3 = ~dec_12[7] & clk;

  always @(posedge clk3) begin
    p0_0_G4_mul0_G16_mul0_G256_inv0_reg3 <= t1_a0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk4;
  assign clk4 = ~dec_12[7] & clk;

  always @(posedge clk4) begin
    p0_0_G4_mul0_G16_mul0_G256_inv0_reg4 <= t12_c0_G4_mul0_G16_mul0_G256_inv0;
  end

  assign t27_a0_G16_mul0_G256_inv0 = a0_0_G16_mul0_G256_inv0 >> dec_2_inp;
  assign t28_b0_G16_mul0_G256_inv0 = ~(~a0_G256_inv0 | ~dec_3_inp);
  assign t26_axorb_0_G16_mul0_G256_inv0 = t27_a0_G16_mul0_G256_inv0 ^ t28_b0_G16_mul0_G256_inv0;
  assign t29_dec_2_inp = dec_2;
  assign t25_a0_0_G4_mul0_G16_mul0_G256_inv0 = t26_axorb_0_G16_mul0_G256_inv0 & t29_dec_2_inp;
  assign t30_dec_1_inp = dec_1;
  assign t24_a0_G4_mul0_G16_mul0_G256_inv0 = ~(~(t25_a0_0_G4_mul0_G16_mul0_G256_inv0 >> t30_dec_1_inp));
  assign t34_a0_0_G16_mul0_G256_inv0 = ~(~a0_G256_inv0 | ~dec_12_inp);
  assign t35_dec_2_inp = dec_2;
  assign t33_a0_G16_mul0_G256_inv0 = ~(~(t34_a0_0_G16_mul0_G256_inv0 >> t35_dec_2_inp));
  assign t37_a0_G256_inv0 = a0_0_G256_inv0 >> dec_4_inp;
  assign t38_dec_3_inp = ~(~dec_3);
  assign t36_b0_G16_mul0_G256_inv0 = ~(~t37_a0_G256_inv0 | ~t38_dec_3_inp);
  assign t32_axorb_0_G16_mul0_G256_inv0 = t33_a0_G16_mul0_G256_inv0 ^ t36_b0_G16_mul0_G256_inv0;
  assign t39_dec_1_inp = dec_1;
  assign t31_b0_G4_mul0_G16_mul0_G256_inv0 = t32_axorb_0_G16_mul0_G256_inv0 & t39_dec_1_inp;
  assign t23_axorb_0_G4_mul0_G16_mul0_G256_inv0 = t24_a0_G4_mul0_G16_mul0_G256_inv0 ^ ~t31_b0_G4_mul0_G16_mul0_G256_inv0;
  assign t44_c0_G16_mul0_G256_inv0 = c0_0_G16_mul0_G256_inv0 >> dec_2_inp;
  assign t45_d0_G16_mul0_G256_inv0 = ~(~b0_G256_inv0 | ~dec_3_inp);
  assign t43_cxord_0_G16_mul0_G256_inv0 = ~(t44_c0_G16_mul0_G256_inv0 ^ ~t45_d0_G16_mul0_G256_inv0);
  assign t46_dec_2_inp = dec_2;
  assign t42_c0_0_G4_mul0_G16_mul0_G256_inv0 = ~(~t43_cxord_0_G16_mul0_G256_inv0 | ~t46_dec_2_inp);
  assign t47_dec_1_inp = ~(~dec_1);
  assign t41_c0_G4_mul0_G16_mul0_G256_inv0 = ~(~(t42_c0_0_G4_mul0_G16_mul0_G256_inv0 >> t47_dec_1_inp));
  assign t51_c0_0_G16_mul0_G256_inv0 = ~(~b0_G256_inv0 | ~dec_12_inp);
  assign t52_dec_2_inp = ~(~dec_2);
  assign t50_c0_G16_mul0_G256_inv0 = ~(~(t51_c0_0_G16_mul0_G256_inv0 >> t52_dec_2_inp));
  assign t54_b0_G256_inv0 = ~(~t2 | ~dec_15_inp);
  assign t55_dec_3_inp = dec_3;
  assign t53_d0_G16_mul0_G256_inv0 = t54_b0_G256_inv0 & t55_dec_3_inp;
  assign t49_cxord_0_G16_mul0_G256_inv0 = ~(~t50_c0_G16_mul0_G256_inv0 ^ t53_d0_G16_mul0_G256_inv0);
  assign t56_dec_1_inp = ~(~dec_1);
  assign t48_d0_G4_mul0_G16_mul0_G256_inv0 = t49_cxord_0_G16_mul0_G256_inv0 & t56_dec_1_inp;
  assign t40_cxord_0_G4_mul0_G16_mul0_G256_inv0 = t41_c0_G4_mul0_G16_mul0_G256_inv0 ^ ~t48_d0_G4_mul0_G16_mul0_G256_inv0;
  wire clk5;
  assign clk5 = dec_243[2] & clk;

  always @(posedge clk5) begin
    e0_G4_mul0_G16_mul0_G256_inv0_reg5 <= axorb_0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk6;
  assign clk6 = dec_243[2] & clk;

  always @(posedge clk6) begin
    e0_G4_mul0_G16_mul0_G256_inv0_reg6 <= cxord_0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk7;
  assign clk7 = ~dec_243[2] & clk;

  always @(posedge clk7) begin
    e0_G4_mul0_G16_mul0_G256_inv0_reg7 <= t23_axorb_0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk8;
  assign clk8 = ~dec_243[2] & clk;

  always @(posedge clk8) begin
    e0_G4_mul0_G16_mul0_G256_inv0_reg8 <= t40_cxord_0_G4_mul0_G16_mul0_G256_inv0;
  end

  assign t61_a0_G256_inv0 = ~(~(a0_0_G256_inv0 >> dec_4_inp));
  assign t62_dec_12_inp = dec_12;
  assign t60_a0_0_G16_mul0_G256_inv0 = ~(~t61_a0_G256_inv0 | ~t62_dec_12_inp);
  assign t63_dec_2_inp = ~(~dec_2);
  assign t59_a0_G16_mul0_G256_inv0 = ~(~(t60_a0_0_G16_mul0_G256_inv0 >> t63_dec_2_inp));
  assign t66_a0_0_G256_inv0 = ~(~t2 | ~dec_240_inp);
  assign t67_dec_4_inp = dec_4;
  assign t65_a0_G256_inv0 = ~(~(t66_a0_0_G256_inv0 >> t67_dec_4_inp));
  assign t68_dec_3_inp = dec_3;
  assign t64_b0_G16_mul0_G256_inv0 = t65_a0_G256_inv0 & t68_dec_3_inp;
  assign t58_axorb_0_G16_mul0_G256_inv0 = ~(~t59_a0_G16_mul0_G256_inv0 ^ t64_b0_G16_mul0_G256_inv0);
  assign t69_dec_1_inp = dec_1;
  assign t57_b0_G4_mul0_G16_mul0_G256_inv0 = ~t58_axorb_0_G16_mul0_G256_inv0 | ~t69_dec_1_inp;
  assign t74_b0_G256_inv0 = ~(~t2 | ~dec_15_inp);
  assign t75_dec_12_inp = ~(~dec_12);
  assign t73_c0_0_G16_mul0_G256_inv0 = t74_b0_G256_inv0 & t75_dec_12_inp;
  assign t76_dec_2_inp = dec_2;
  assign t72_c0_G16_mul0_G256_inv0 = t73_c0_0_G16_mul0_G256_inv0 >> t76_dec_2_inp;
  assign t80_y8_G256_newbasis0 = ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0;
  assign t79_t2 = ~(~t80_y8_G256_newbasis0);
  assign t81_dec_15_inp = ~(~dec_15);
  assign t78_b0_G256_inv0 = ~(~t79_t2 | ~t81_dec_15_inp);
  assign t82_dec_3_inp = dec_3;
  assign t77_d0_G16_mul0_G256_inv0 = t78_b0_G256_inv0 & t82_dec_3_inp;
  assign t71_cxord_0_G16_mul0_G256_inv0 = t72_c0_G16_mul0_G256_inv0 ^ t77_d0_G16_mul0_G256_inv0;
  assign t83_dec_1_inp = dec_1;
  assign t70_d0_G4_mul0_G16_mul0_G256_inv0 = ~t71_cxord_0_G16_mul0_G256_inv0 | ~t83_dec_1_inp;
  wire clk9;
  assign clk9 = dec_152[0] & clk;

  always @(posedge clk9) begin
    q0_0_G4_mul0_G16_mul0_G256_inv0_reg9 <= b0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk10;
  assign clk10 = dec_152[0] & clk;

  always @(posedge clk10) begin
    q0_0_G4_mul0_G16_mul0_G256_inv0_reg10 <= d0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk11;
  assign clk11 = ~dec_152[0] & clk;

  always @(posedge clk11) begin
    q0_0_G4_mul0_G16_mul0_G256_inv0_reg11 <= t57_b0_G4_mul0_G16_mul0_G256_inv0;
  end

  wire clk12;
  assign clk12 = ~dec_152[0] & clk;

  always @(posedge clk12) begin
    q0_0_G4_mul0_G16_mul0_G256_inv0_reg12 <= t70_d0_G4_mul0_G16_mul0_G256_inv0;
  end

  assign t88_a0_G256_inv0 = a0_0_G256_inv0 >> dec_4_inp;
  assign t89_dec_12_inp = ~(~dec_12);
  assign t87_a0_0_G16_mul0_G256_inv0 = t88_a0_G256_inv0 & t89_dec_12_inp;
  assign t90_dec_2_inp = ~(~dec_2);
  assign t86_a0_G16_mul0_G256_inv0 = t87_a0_0_G16_mul0_G256_inv0 >> t90_dec_2_inp;
  assign t91_dec_2_inp = ~(~dec_2);
  assign t85_a0_0_G4_mul1_G16_mul0_G256_inv0 = ~(~t86_a0_G16_mul0_G256_inv0 | ~t91_dec_2_inp);
  assign t92_dec_1_inp = ~(~dec_1);
  assign t84_a0_G4_mul1_G16_mul0_G256_inv0 = ~(t85_a0_0_G4_mul1_G16_mul0_G256_inv0 >> t92_dec_1_inp);
  assign t97_b0_G256_inv0 = ~(~t2 | ~dec_15_inp);
  assign t98_dec_12_inp = dec_12;
  assign t96_c0_0_G16_mul0_G256_inv0 = t97_b0_G256_inv0 & t98_dec_12_inp;
  assign t99_dec_2_inp = dec_2;
  assign t95_c0_G16_mul0_G256_inv0 = ~(~(t96_c0_0_G16_mul0_G256_inv0 >> t99_dec_2_inp));
  assign t100_dec_2_inp = dec_2;
  assign t94_c0_0_G4_mul1_G16_mul0_G256_inv0 = ~(~t95_c0_G16_mul0_G256_inv0 | ~t100_dec_2_inp);
  assign t101_dec_1_inp = dec_1;
  assign t93_c0_G4_mul1_G16_mul0_G256_inv0 = ~(t94_c0_0_G4_mul1_G16_mul0_G256_inv0 >> t101_dec_1_inp);
  wire clk13;
  assign clk13 = dec_243[5] & clk;

  always @(posedge clk13) begin
    p0_0_G4_mul1_G16_mul0_G256_inv0_reg13 <= a0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk14;
  assign clk14 = dec_243[5] & clk;

  always @(posedge clk14) begin
    p0_0_G4_mul1_G16_mul0_G256_inv0_reg14 <= c0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk15;
  assign clk15 = ~dec_243[5] & clk;

  always @(posedge clk15) begin
    p0_0_G4_mul1_G16_mul0_G256_inv0_reg15 <= t84_a0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk16;
  assign clk16 = ~dec_243[5] & clk;

  always @(posedge clk16) begin
    p0_0_G4_mul1_G16_mul0_G256_inv0_reg16 <= t93_c0_G4_mul1_G16_mul0_G256_inv0;
  end

  assign t106_a0_0_G16_mul0_G256_inv0 = a0_G256_inv0 & dec_12_inp;
  assign t107_dec_2_inp = dec_2;
  assign t105_a0_G16_mul0_G256_inv0 = t106_a0_0_G16_mul0_G256_inv0 >> t107_dec_2_inp;
  assign t108_dec_2_inp = dec_2;
  assign t104_a0_0_G4_mul1_G16_mul0_G256_inv0 = ~(~t105_a0_G16_mul0_G256_inv0 | ~t108_dec_2_inp);
  assign t109_dec_1_inp = ~(~dec_1);
  assign t103_a0_G4_mul1_G16_mul0_G256_inv0 = t104_a0_0_G4_mul1_G16_mul0_G256_inv0 >> t109_dec_1_inp;
  assign t113_a0_G256_inv0 = a0_0_G256_inv0 >> dec_4_inp;
  assign t114_dec_12_inp = dec_12;
  assign t112_a0_0_G16_mul0_G256_inv0 = ~(~t113_a0_G256_inv0 | ~t114_dec_12_inp);
  assign t115_dec_2_inp = dec_2;
  assign t111_a0_G16_mul0_G256_inv0 = t112_a0_0_G16_mul0_G256_inv0 >> t115_dec_2_inp;
  assign t116_dec_1_inp = dec_1;
  assign t110_b0_G4_mul1_G16_mul0_G256_inv0 = ~(~t111_a0_G16_mul0_G256_inv0 | ~t116_dec_1_inp);
  assign t102_axorb_0_G4_mul1_G16_mul0_G256_inv0 = ~(~(~t103_a0_G4_mul1_G16_mul0_G256_inv0)) ^ t110_b0_G4_mul1_G16_mul0_G256_inv0;
  assign t121_c0_0_G16_mul0_G256_inv0 = ~(~b0_G256_inv0 | ~dec_12_inp);
  assign t122_dec_2_inp = dec_2;
  assign t120_c0_G16_mul0_G256_inv0 = t121_c0_0_G16_mul0_G256_inv0 >> t122_dec_2_inp;
  assign t123_dec_2_inp = dec_2;
  assign t119_c0_0_G4_mul1_G16_mul0_G256_inv0 = ~(~t120_c0_G16_mul0_G256_inv0 | ~t123_dec_2_inp);
  assign t124_dec_1_inp = dec_1;
  assign t118_c0_G4_mul1_G16_mul0_G256_inv0 = ~(~(t119_c0_0_G4_mul1_G16_mul0_G256_inv0 >> t124_dec_1_inp));
  assign t128_b0_G256_inv0 = ~(~t2 | ~dec_15_inp);
  assign t129_dec_12_inp = ~(~dec_12);
  assign t127_c0_0_G16_mul0_G256_inv0 = t128_b0_G256_inv0 & t129_dec_12_inp;
  assign t130_dec_2_inp = ~(~dec_2);
  assign t126_c0_G16_mul0_G256_inv0 = ~(~(t127_c0_0_G16_mul0_G256_inv0 >> t130_dec_2_inp));
  assign t131_dec_1_inp = ~(~dec_1);
  assign t125_d0_G4_mul1_G16_mul0_G256_inv0 = ~(~t126_c0_G16_mul0_G256_inv0 | ~t131_dec_1_inp);
  assign t117_cxord_0_G4_mul1_G16_mul0_G256_inv0 = ~(~t118_c0_G4_mul1_G16_mul0_G256_inv0) ^ ~t125_d0_G4_mul1_G16_mul0_G256_inv0;
  wire clk17;
  assign clk17 = dec_9[7] & clk;

  always @(posedge clk17) begin
    e0_G4_mul1_G16_mul0_G256_inv0_reg17 <= a0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk18;
  assign clk18 = dec_9[7] & clk;

  always @(posedge clk18) begin
    e0_G4_mul1_G16_mul0_G256_inv0_reg18 <= b0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk19;
  assign clk19 = dec_9[7] & clk;

  always @(posedge clk19) begin
    e0_G4_mul1_G16_mul0_G256_inv0_reg19 <= c0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk20;
  assign clk20 = dec_9[7] & clk;

  always @(posedge clk20) begin
    e0_G4_mul1_G16_mul0_G256_inv0_reg20 <= d0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk21;
  assign clk21 = ~dec_9[7] & clk;

  always @(posedge clk21) begin
    e0_G4_mul1_G16_mul0_G256_inv0_reg21 <= t102_axorb_0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk22;
  assign clk22 = ~dec_9[7] & clk;

  always @(posedge clk22) begin
    e0_G4_mul1_G16_mul0_G256_inv0_reg22 <= t117_cxord_0_G4_mul1_G16_mul0_G256_inv0;
  end

  assign t136_a0_0_G256_inv0 = t2 & dec_240_inp;
  assign t137_dec_4_inp = dec_4;
  assign t135_a0_G256_inv0 = ~(~(t136_a0_0_G256_inv0 >> t137_dec_4_inp));
  assign t138_dec_12_inp = dec_12;
  assign t134_a0_0_G16_mul0_G256_inv0 = ~(~t135_a0_G256_inv0 | ~t138_dec_12_inp);
  assign t139_dec_2_inp = ~(~dec_2);
  assign t133_a0_G16_mul0_G256_inv0 = t134_a0_0_G16_mul0_G256_inv0 >> t139_dec_2_inp;
  assign t140_dec_1_inp = ~(~dec_1);
  assign t132_b0_G4_mul1_G16_mul0_G256_inv0 = ~t133_a0_G16_mul0_G256_inv0 | ~t140_dec_1_inp;
  assign t146_y8_G256_newbasis0 = ~(~ny8_G256_newbasis0 + (~tempyIntoNegCond8_G256_newbasis0 + 1));
  assign t145_t2 = t146_y8_G256_newbasis0;
  assign t147_dec_15_inp = dec_15;
  assign t144_b0_G256_inv0 = t145_t2 & t147_dec_15_inp;
  assign t148_dec_12_inp = ~(~dec_12);
  assign t143_c0_0_G16_mul0_G256_inv0 = ~(~t144_b0_G256_inv0 | ~t148_dec_12_inp);
  assign t149_dec_2_inp = ~(~dec_2);
  assign t142_c0_G16_mul0_G256_inv0 = t143_c0_0_G16_mul0_G256_inv0 >> t149_dec_2_inp;
  assign t150_dec_1_inp = dec_1;
  assign t141_d0_G4_mul1_G16_mul0_G256_inv0 = ~t142_c0_G16_mul0_G256_inv0 | ~t150_dec_1_inp;
  wire clk23;
  assign clk23 = dec_243[6] & clk;

  always @(posedge clk23) begin
    q0_0_G4_mul1_G16_mul0_G256_inv0_reg23 <= b0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk24;
  assign clk24 = dec_243[6] & clk;

  always @(posedge clk24) begin
    q0_0_G4_mul1_G16_mul0_G256_inv0_reg24 <= d0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk25;
  assign clk25 = ~dec_243[6] & clk;

  always @(posedge clk25) begin
    q0_0_G4_mul1_G16_mul0_G256_inv0_reg25 <= t132_b0_G4_mul1_G16_mul0_G256_inv0;
  end

  wire clk26;
  assign clk26 = ~dec_243[6] & clk;

  always @(posedge clk26) begin
    q0_0_G4_mul1_G16_mul0_G256_inv0_reg26 <= t141_d0_G4_mul1_G16_mul0_G256_inv0;
  end

  assign t155_a0_0_G256_inv0 = t2 & dec_240_inp;
  assign t156_dec_4_inp = ~(~dec_4);
  assign t154_a0_G256_inv0 = t155_a0_0_G256_inv0 >> t156_dec_4_inp;
  assign t157_dec_3_inp = ~(~dec_3);
  assign t153_b0_G16_mul0_G256_inv0 = t154_a0_G256_inv0 & t157_dec_3_inp;
  assign t158_dec_2_inp = dec_2;
  assign t152_a0_0_G4_mul2_G16_mul0_G256_inv0 = t153_b0_G16_mul0_G256_inv0 & t158_dec_2_inp;
  assign t159_dec_1_inp = ~(~dec_1);
  assign t151_a0_G4_mul2_G16_mul0_G256_inv0 = ~(~(t152_a0_0_G4_mul2_G16_mul0_G256_inv0 >> t159_dec_1_inp));
  assign t165_y8_G256_newbasis0 = ~(~ny8_G256_newbasis0 + (~tempyIntoNegCond8_G256_newbasis0 + 1));
  assign t164_t2 = t165_y8_G256_newbasis0;
  assign t166_dec_15_inp = dec_15;
  assign t163_b0_G256_inv0 = t164_t2 & t166_dec_15_inp;
  assign t167_dec_3_inp = ~(~dec_3);
  assign t162_d0_G16_mul0_G256_inv0 = t163_b0_G256_inv0 & t167_dec_3_inp;
  assign t168_dec_2_inp = ~(~dec_2);
  assign t161_c0_0_G4_mul2_G16_mul0_G256_inv0 = ~(~t162_d0_G16_mul0_G256_inv0 | ~t168_dec_2_inp);
  assign t169_dec_1_inp = ~(~dec_1);
  assign t160_c0_G4_mul2_G16_mul0_G256_inv0 = t161_c0_0_G4_mul2_G16_mul0_G256_inv0 >> t169_dec_1_inp;
  wire clk27;
  assign clk27 = dec_12[0] & clk;

  always @(posedge clk27) begin
    p0_0_G4_mul2_G16_mul0_G256_inv0_reg27 <= a0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk28;
  assign clk28 = dec_12[0] & clk;

  always @(posedge clk28) begin
    p0_0_G4_mul2_G16_mul0_G256_inv0_reg28 <= c0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk29;
  assign clk29 = ~dec_12[0] & clk;

  always @(posedge clk29) begin
    p0_0_G4_mul2_G16_mul0_G256_inv0_reg29 <= t151_a0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk30;
  assign clk30 = ~dec_12[0] & clk;

  always @(posedge clk30) begin
    p0_0_G4_mul2_G16_mul0_G256_inv0_reg30 <= t160_c0_G4_mul2_G16_mul0_G256_inv0;
  end

  assign t174_a0_G256_inv0 = ~(~(a0_0_G256_inv0 >> dec_4_inp));
  assign t175_dec_3_inp = ~(~dec_3);
  assign t173_b0_G16_mul0_G256_inv0 = ~(~t174_a0_G256_inv0 | ~t175_dec_3_inp);
  assign t176_dec_2_inp = dec_2;
  assign t172_a0_0_G4_mul2_G16_mul0_G256_inv0 = t173_b0_G16_mul0_G256_inv0 & t176_dec_2_inp;
  assign t177_dec_1_inp = ~(~dec_1);
  assign t171_a0_G4_mul2_G16_mul0_G256_inv0 = ~(t172_a0_0_G4_mul2_G16_mul0_G256_inv0 >> t177_dec_1_inp);
  assign t181_a0_0_G256_inv0 = t2 & dec_240_inp;
  assign t182_dec_4_inp = dec_4;
  assign t180_a0_G256_inv0 = t181_a0_0_G256_inv0 >> t182_dec_4_inp;
  assign t183_dec_3_inp = ~(~dec_3);
  assign t179_b0_G16_mul0_G256_inv0 = ~(~t180_a0_G256_inv0 | ~t183_dec_3_inp);
  assign t184_dec_1_inp = ~(~dec_1);
  assign t178_b0_G4_mul2_G16_mul0_G256_inv0 = t179_b0_G16_mul0_G256_inv0 & t184_dec_1_inp;
  assign t170_axorb_0_G4_mul2_G16_mul0_G256_inv0 = ~(~t171_a0_G4_mul2_G16_mul0_G256_inv0) ^ t178_b0_G4_mul2_G16_mul0_G256_inv0;
  assign t189_b0_G256_inv0 = t2 & dec_15_inp;
  assign t190_dec_3_inp = dec_3;
  assign t188_d0_G16_mul0_G256_inv0 = t189_b0_G256_inv0 & t190_dec_3_inp;
  assign t191_dec_2_inp = ~(~dec_2);
  assign t187_c0_0_G4_mul2_G16_mul0_G256_inv0 = ~(~t188_d0_G16_mul0_G256_inv0 | ~t191_dec_2_inp);
  assign t192_dec_1_inp = ~(~dec_1);
  assign t186_c0_G4_mul2_G16_mul0_G256_inv0 = ~(t187_c0_0_G4_mul2_G16_mul0_G256_inv0 >> t192_dec_1_inp);
  assign t197_y8_G256_newbasis0 = ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0;
  assign t196_t2 = ~(~t197_y8_G256_newbasis0);
  assign t198_dec_15_inp = dec_15;
  assign t195_b0_G256_inv0 = ~(~t196_t2 | ~t198_dec_15_inp);
  assign t199_dec_3_inp = dec_3;
  assign t194_d0_G16_mul0_G256_inv0 = ~(~t195_b0_G256_inv0 | ~t199_dec_3_inp);
  assign t200_dec_1_inp = dec_1;
  assign t193_d0_G4_mul2_G16_mul0_G256_inv0 = t194_d0_G16_mul0_G256_inv0 & t200_dec_1_inp;
  assign t185_cxord_0_G4_mul2_G16_mul0_G256_inv0 = ~t186_c0_G4_mul2_G16_mul0_G256_inv0 ^ ~t193_d0_G4_mul2_G16_mul0_G256_inv0;
  wire clk31;
  assign clk31 = dec_0[5] & clk;

  always @(posedge clk31) begin
    e0_G4_mul2_G16_mul0_G256_inv0_reg31 <= a0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk32;
  assign clk32 = dec_0[5] & clk;

  always @(posedge clk32) begin
    e0_G4_mul2_G16_mul0_G256_inv0_reg32 <= b0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk33;
  assign clk33 = dec_0[5] & clk;

  always @(posedge clk33) begin
    e0_G4_mul2_G16_mul0_G256_inv0_reg33 <= c0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk34;
  assign clk34 = dec_0[5] & clk;

  always @(posedge clk34) begin
    e0_G4_mul2_G16_mul0_G256_inv0_reg34 <= d0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk35;
  assign clk35 = ~dec_0[5] & clk;

  always @(posedge clk35) begin
    e0_G4_mul2_G16_mul0_G256_inv0_reg35 <= t170_axorb_0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk36;
  assign clk36 = ~dec_0[5] & clk;

  always @(posedge clk36) begin
    e0_G4_mul2_G16_mul0_G256_inv0_reg36 <= t185_cxord_0_G4_mul2_G16_mul0_G256_inv0;
  end

  assign t206_y8_G256_newbasis0 = ~(~ny8_G256_newbasis0 + (~tempyIntoNegCond8_G256_newbasis0 + 1));
  assign t205_t2 = ~(~t206_y8_G256_newbasis0);
  assign t207_dec_240_inp = dec_240;
  assign t204_a0_0_G256_inv0 = t205_t2 & t207_dec_240_inp;
  assign t208_dec_4_inp = dec_4;
  assign t203_a0_G256_inv0 = t204_a0_0_G256_inv0 >> t208_dec_4_inp;
  assign t209_dec_3_inp = dec_3;
  assign t202_b0_G16_mul0_G256_inv0 = ~(~t203_a0_G256_inv0 | ~t209_dec_3_inp);
  assign t210_dec_1_inp = ~(~dec_1);
  assign t201_b0_G4_mul2_G16_mul0_G256_inv0 = ~t202_b0_G16_mul0_G256_inv0 | ~t210_dec_1_inp;
  assign t216_ny8_G256_newbasis0 = cond8_G256_newbasis0 * yxorb8_G256_newbasis0;
  assign t217_tempyIntoNegCond8_G256_newbasis0 = tempy8_G256_newbasis0 * negCond8_G256_newbasis0;
  assign t215_y8_G256_newbasis0 = ~(~t216_ny8_G256_newbasis0 + (~t217_tempyIntoNegCond8_G256_newbasis0 + 1));
  assign t214_t2 = ~(~t215_y8_G256_newbasis0);
  assign t218_dec_15_inp = dec_15;
  assign t213_b0_G256_inv0 = t214_t2 & t218_dec_15_inp;
  assign t219_dec_3_inp = ~(~dec_3);
  assign t212_d0_G16_mul0_G256_inv0 = t213_b0_G256_inv0 & t219_dec_3_inp;
  assign t220_dec_1_inp = ~(~dec_1);
  assign t211_d0_G4_mul2_G16_mul0_G256_inv0 = ~t212_d0_G16_mul0_G256_inv0 | ~t220_dec_1_inp;
  wire clk37;
  assign clk37 = dec_169[1] & clk;

  always @(posedge clk37) begin
    q0_0_G4_mul2_G16_mul0_G256_inv0_reg37 <= b0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk38;
  assign clk38 = dec_169[1] & clk;

  always @(posedge clk38) begin
    q0_0_G4_mul2_G16_mul0_G256_inv0_reg38 <= d0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk39;
  assign clk39 = ~dec_169[1] & clk;

  always @(posedge clk39) begin
    q0_0_G4_mul2_G16_mul0_G256_inv0_reg39 <= t201_b0_G4_mul2_G16_mul0_G256_inv0;
  end

  wire clk40;
  assign clk40 = ~dec_169[1] & clk;

  always @(posedge clk40) begin
    q0_0_G4_mul2_G16_mul0_G256_inv0_reg40 <= t211_d0_G4_mul2_G16_mul0_G256_inv0;
  end

  assign t225_c0xord0_G256_inv0 = ~(y_reg141 ^ ~d0_G256_inv0);
  assign t226_dec_12_inp = ~(~dec_12);
  assign t224_a0_0_G16_inv0_G256_inv0 = ~(~t225_c0xord0_G256_inv0 | y_reg142);
  assign t227_dec_2_inp = ~(~dec_2);
  assign t223_a0_G16_inv0_G256_inv0 = t224_a0_0_G16_inv0_G256_inv0 >> y_reg143;
  assign t228_dec_2_inp = dec_2;
  assign t222_a0_0_G4_mul3_G16_inv0_G256_inv0 = ~(~t223_a0_G16_inv0_G256_inv0 | y_reg144);
  assign t229_dec_1_inp = dec_1;
  assign t221_a0_G4_mul3_G16_inv0_G256_inv0 = ~(~(t222_a0_0_G4_mul3_G16_inv0_G256_inv0 >> y_reg145));
  assign t234_c0_G256_inv0 = p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0;
  assign t235_d0_G256_inv0 = p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0;
  assign t233_c0xord0_G256_inv0 = y_reg146 ^ t235_d0_G256_inv0;
  assign t236_dec_3_inp = dec_3;
  assign t232_b0_G16_inv0_G256_inv0 = t233_c0xord0_G256_inv0 & y_reg147;
  assign t237_dec_2_inp = ~(~dec_2);
  assign t231_c0_0_G4_mul3_G16_inv0_G256_inv0 = t232_b0_G16_inv0_G256_inv0 & y_reg148;
  assign t238_dec_1_inp = ~(~dec_1);
  assign t230_c0_G4_mul3_G16_inv0_G256_inv0 = ~(~(t231_c0_0_G4_mul3_G16_inv0_G256_inv0 >> y_reg149));
  wire clk41;
  assign clk41 = dec_36[5] & clk;

  always @(posedge clk41) begin
    p0_0_G4_mul3_G16_inv0_G256_inv0_reg41 <= a0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk42;
  assign clk42 = dec_36[5] & clk;

  always @(posedge clk42) begin
    p0_0_G4_mul3_G16_inv0_G256_inv0_reg42 <= c0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk43;
  assign clk43 = ~dec_36[5] & clk;

  always @(posedge clk43) begin
    p0_0_G4_mul3_G16_inv0_G256_inv0_reg43 <= t221_a0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk44;
  assign clk44 = ~dec_36[5] & clk;

  always @(posedge clk44) begin
    p0_0_G4_mul3_G16_inv0_G256_inv0_reg44 <= t230_c0_G4_mul3_G16_inv0_G256_inv0;
  end

  assign t243_a0_0_G16_inv0_G256_inv0 = ~(~c0xord0_G256_inv0 | y_reg154);
  assign t244_dec_2_inp = ~(~dec_2);
  assign t242_a0_G16_inv0_G256_inv0 = ~(~(t243_a0_0_G16_inv0_G256_inv0 >> y_reg155));
  assign t245_dec_2_inp = dec_2;
  assign t241_a0_0_G4_mul3_G16_inv0_G256_inv0 = ~(~t242_a0_G16_inv0_G256_inv0 | y_reg156);
  assign t246_dec_1_inp = dec_1;
  assign t240_a0_G4_mul3_G16_inv0_G256_inv0 = ~(~(t241_a0_0_G4_mul3_G16_inv0_G256_inv0 >> y_reg157));
  assign t250_c0xord0_G256_inv0 = y_reg158 ^ d0_G256_inv0;
  assign t251_dec_12_inp = dec_12;
  assign t249_a0_0_G16_inv0_G256_inv0 = t250_c0xord0_G256_inv0 & y_reg159;
  assign t252_dec_2_inp = dec_2;
  assign t248_a0_G16_inv0_G256_inv0 = ~(~(t249_a0_0_G16_inv0_G256_inv0 >> y_reg160));
  assign t253_dec_1_inp = ~(~dec_1);
  assign t247_b0_G4_mul3_G16_inv0_G256_inv0 = ~(~t248_a0_G16_inv0_G256_inv0 | y_reg161);
  assign t239_axorb_0_G4_mul3_G16_inv0_G256_inv0 = ~(~t240_a0_G4_mul3_G16_inv0_G256_inv0 ^ t247_b0_G4_mul3_G16_inv0_G256_inv0);
  assign t258_c0xord0_G256_inv0 = y_reg162 ^ d0_G256_inv0;
  assign t259_dec_3_inp = dec_3;
  assign t257_b0_G16_inv0_G256_inv0 = ~(~t258_c0xord0_G256_inv0 | y_reg163);
  assign t260_dec_2_inp = ~(~dec_2);
  assign t256_c0_0_G4_mul3_G16_inv0_G256_inv0 = ~(~t257_b0_G16_inv0_G256_inv0 | y_reg164);
  assign t261_dec_1_inp = ~(~dec_1);
  assign t255_c0_G4_mul3_G16_inv0_G256_inv0 = t256_c0_0_G4_mul3_G16_inv0_G256_inv0 >> y_reg165;
  assign t265_c0_G256_inv0 = ~(~p0ls2_G16_sq_scl0_G256_inv0 & ~q0_G16_sq_scl0_G256_inv0);
  assign t266_d0_G256_inv0 = ~(~p0ls2_G16_mul0_G256_inv0 & ~q0_G16_mul0_G256_inv0);
  assign t264_c0xord0_G256_inv0 = y_reg166 ^ t266_d0_G256_inv0;
  assign t267_dec_3_inp = dec_3;
  assign t263_b0_G16_inv0_G256_inv0 = t264_c0xord0_G256_inv0 & y_reg167;
  assign t268_dec_1_inp = dec_1;
  assign t262_d0_G4_mul3_G16_inv0_G256_inv0 = t263_b0_G16_inv0_G256_inv0 & y_reg168;
  assign t254_cxord_0_G4_mul3_G16_inv0_G256_inv0 = t255_c0_G4_mul3_G16_inv0_G256_inv0 ^ t262_d0_G4_mul3_G16_inv0_G256_inv0;
  wire clk45;
  assign clk45 = r[13] & clk;

  always @(posedge clk45) begin
    e0_G4_mul3_G16_inv0_G256_inv0_reg45 <= a0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk46;
  assign clk46 = r[13] & clk;

  always @(posedge clk46) begin
    e0_G4_mul3_G16_inv0_G256_inv0_reg46 <= b0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk47;
  assign clk47 = r[13] & clk;

  always @(posedge clk47) begin
    e0_G4_mul3_G16_inv0_G256_inv0_reg47 <= c0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk48;
  assign clk48 = r[13] & clk;

  always @(posedge clk48) begin
    e0_G4_mul3_G16_inv0_G256_inv0_reg48 <= d0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk49;
  assign clk49 = ~r[13] & clk;

  always @(posedge clk49) begin
    e0_G4_mul3_G16_inv0_G256_inv0_reg49 <= t239_axorb_0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk50;
  assign clk50 = ~r[13] & clk;

  always @(posedge clk50) begin
    e0_G4_mul3_G16_inv0_G256_inv0_reg50 <= t254_cxord_0_G4_mul3_G16_inv0_G256_inv0;
  end

  assign t273_c0_G256_inv0 = ~(~p0ls2_G16_sq_scl0_G256_inv0 & ~q0_G16_sq_scl0_G256_inv0);
  assign t274_d0_G256_inv0 = p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0;
  assign t272_c0xord0_G256_inv0 = y_reg173 ^ t274_d0_G256_inv0;
  assign t275_dec_12_inp = ~(~dec_12);
  assign t271_a0_0_G16_inv0_G256_inv0 = ~(~t272_c0xord0_G256_inv0 | y_reg174);
  assign t276_dec_2_inp = dec_2;
  assign t270_a0_G16_inv0_G256_inv0 = t271_a0_0_G16_inv0_G256_inv0 >> y_reg175;
  assign t277_dec_1_inp = dec_1;
  assign t269_b0_G4_mul3_G16_inv0_G256_inv0 = ~t270_a0_G16_inv0_G256_inv0 | y_reg176;
  assign t282_p0ls2_G16_sq_scl0_G256_inv0 = p0_G16_sq_scl0_G256_inv0 << dec_2_inp;
  assign t283_q0_G16_sq_scl0_G256_inv0 = ~(~p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 & ~q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
  assign t281_c0_G256_inv0 = ~(~t282_p0ls2_G16_sq_scl0_G256_inv0 & ~t283_q0_G16_sq_scl0_G256_inv0);
  assign t285_p0ls2_G16_mul0_G256_inv0 = ~(~(p0_G16_mul0_G256_inv0 << y_reg177));
  assign t286_q0_G16_mul0_G256_inv0 = ~(~q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
  assign t284_d0_G256_inv0 = t285_p0ls2_G16_mul0_G256_inv0 | t286_q0_G16_mul0_G256_inv0;
  assign t280_c0xord0_G256_inv0 = y_reg178 ^ t284_d0_G256_inv0;
  assign t287_dec_3_inp = ~(~dec_3);
  assign t279_b0_G16_inv0_G256_inv0 = ~t280_c0xord0_G256_inv0 | y_reg179;
  assign t288_dec_1_inp = ~dec_1;
  assign t278_d0_G4_mul3_G16_inv0_G256_inv0 = t279_b0_G16_inv0_G256_inv0 | y_reg180;
  wire clk51;
  assign clk51 = dec_242[4] & clk;

  always @(posedge clk51) begin
    q0_0_G4_mul3_G16_inv0_G256_inv0_reg51 <= b0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk52;
  assign clk52 = dec_242[4] & clk;

  always @(posedge clk52) begin
    q0_0_G4_mul3_G16_inv0_G256_inv0_reg52 <= d0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk53;
  assign clk53 = ~dec_242[4] & clk;

  always @(posedge clk53) begin
    q0_0_G4_mul3_G16_inv0_G256_inv0_reg53 <= t269_b0_G4_mul3_G16_inv0_G256_inv0;
  end

  wire clk54;
  assign clk54 = ~dec_242[4] & clk;

  always @(posedge clk54) begin
    q0_0_G4_mul3_G16_inv0_G256_inv0_reg54 <= t278_d0_G4_mul3_G16_inv0_G256_inv0;
  end

  assign t293_b0_G4_sq3_G16_inv0_G256_inv0 = ~(~c0xord0_G16_inv0_G256_inv0 | y_reg183);
  assign t294_dec_1_inp = ~(~dec_1);
  assign t292_b0ls1_G4_sq3_G16_inv0_G256_inv0 = t293_b0_G4_sq3_G16_inv0_G256_inv0 << y_reg185;
  assign t296_a0_0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg187;
  assign t297_dec_1_inp = ~(~dec_1);
  assign t295_a0_G4_sq3_G16_inv0_G256_inv0 = t296_a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg189;
  assign t291_e0_G16_inv0_G256_inv0 = t292_b0ls1_G4_sq3_G16_inv0_G256_inv0 | t295_a0_G4_sq3_G16_inv0_G256_inv0;
  assign t298_dec_2_inp = dec_2;
  assign t290_a0_0_G4_mul4_G16_inv0_G256_inv0 = ~(~t291_e0_G16_inv0_G256_inv0 | y_reg191);
  assign t299_dec_1_inp = ~(~dec_1);
  assign t289_a0_G4_mul4_G16_inv0_G256_inv0 = ~(t290_a0_0_G4_mul4_G16_inv0_G256_inv0 >> y_reg193);
  assign t304_c0_G256_inv0 = p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0;
  assign t305_d0_G256_inv0 = p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0;
  assign t303_c0xord0_G256_inv0 = ~(y_reg194 ^ t305_d0_G256_inv0);
  assign t306_dec_3_inp = ~(~dec_3);
  assign t302_b0_G16_inv0_G256_inv0 = t303_c0xord0_G256_inv0 & y_reg195;
  assign t307_dec_2_inp = ~(~dec_2);
  assign t301_c0_0_G4_mul4_G16_inv0_G256_inv0 = t302_b0_G16_inv0_G256_inv0 & y_reg196;
  assign t308_dec_1_inp = ~(~dec_1);
  assign t300_c0_G4_mul4_G16_inv0_G256_inv0 = ~(t301_c0_0_G4_mul4_G16_inv0_G256_inv0 >> y_reg197);
  wire clk55;
  assign clk55 = t[4] & clk;

  always @(posedge clk55) begin
    p0_0_G4_mul4_G16_inv0_G256_inv0_reg55 <= a0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk56;
  assign clk56 = t[4] & clk;

  always @(posedge clk56) begin
    p0_0_G4_mul4_G16_inv0_G256_inv0_reg56 <= c0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk57;
  assign clk57 = ~t[4] & clk;

  always @(posedge clk57) begin
    p0_0_G4_mul4_G16_inv0_G256_inv0_reg57 <= t289_a0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk58;
  assign clk58 = ~t[4] & clk;

  always @(posedge clk58) begin
    p0_0_G4_mul4_G16_inv0_G256_inv0_reg58 <= t300_c0_G4_mul4_G16_inv0_G256_inv0;
  end

  assign t313_b0ls1_G4_sq3_G16_inv0_G256_inv0 = b0_G4_sq3_G16_inv0_G256_inv0 << y_reg215;
  assign t314_a0_G4_sq3_G16_inv0_G256_inv0 = a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg217;
  assign t312_e0_G16_inv0_G256_inv0 = t313_b0ls1_G4_sq3_G16_inv0_G256_inv0 | t314_a0_G4_sq3_G16_inv0_G256_inv0;
  assign t315_dec_2_inp = ~(~dec_2);
  assign t311_a0_0_G4_mul4_G16_inv0_G256_inv0 = t312_e0_G16_inv0_G256_inv0 & y_reg219;
  assign t316_dec_1_inp = ~(~dec_1);
  assign t310_a0_G4_mul4_G16_inv0_G256_inv0 = t311_a0_0_G4_mul4_G16_inv0_G256_inv0 >> y_reg221;
  assign t320_b0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg223;
  assign t321_dec_1_inp = ~(~dec_1);
  assign t319_b0ls1_G4_sq3_G16_inv0_G256_inv0 = t320_b0_G4_sq3_G16_inv0_G256_inv0 << y_reg225;
  assign t323_a0_0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg227;
  assign t324_dec_1_inp = dec_1;
  assign t322_a0_G4_sq3_G16_inv0_G256_inv0 = t323_a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg229;
  assign t318_e0_G16_inv0_G256_inv0 = ~(~t319_b0ls1_G4_sq3_G16_inv0_G256_inv0 & ~t322_a0_G4_sq3_G16_inv0_G256_inv0);
  assign t325_dec_1_inp = ~(~dec_1);
  assign t317_b0_G4_mul4_G16_inv0_G256_inv0 = ~(~t318_e0_G16_inv0_G256_inv0 | y_reg231);
  assign t309_axorb_0_G4_mul4_G16_inv0_G256_inv0 = t310_a0_G4_mul4_G16_inv0_G256_inv0 ^ ~t317_b0_G4_mul4_G16_inv0_G256_inv0;
  assign t330_c0xord0_G256_inv0 = ~(y_reg232 ^ d0_G256_inv0);
  assign t331_dec_3_inp = ~(~dec_3);
  assign t329_b0_G16_inv0_G256_inv0 = ~(~t330_c0xord0_G256_inv0 | y_reg233);
  assign t332_dec_2_inp = ~(~dec_2);
  assign t328_c0_0_G4_mul4_G16_inv0_G256_inv0 = ~(~t329_b0_G16_inv0_G256_inv0 | y_reg234);
  assign t333_dec_1_inp = ~(~dec_1);
  assign t327_c0_G4_mul4_G16_inv0_G256_inv0 = ~(~(t328_c0_0_G4_mul4_G16_inv0_G256_inv0 >> y_reg235));
  assign t337_c0_G256_inv0 = ~(~p0ls2_G16_sq_scl0_G256_inv0 & ~q0_G16_sq_scl0_G256_inv0);
  assign t338_d0_G256_inv0 = p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0;
  assign t336_c0xord0_G256_inv0 = ~(y_reg236 ^ t338_d0_G256_inv0);
  assign t339_dec_3_inp = ~(~dec_3);
  assign t335_b0_G16_inv0_G256_inv0 = t336_c0xord0_G256_inv0 & y_reg237;
  assign t340_dec_1_inp = dec_1;
  assign t334_d0_G4_mul4_G16_inv0_G256_inv0 = t335_b0_G16_inv0_G256_inv0 & y_reg238;
  assign t326_cxord_0_G4_mul4_G16_inv0_G256_inv0 = ~t327_c0_G4_mul4_G16_inv0_G256_inv0 ^ t334_d0_G4_mul4_G16_inv0_G256_inv0;
  wire clk59;
  assign clk59 = dec_255[0] & clk;

  always @(posedge clk59) begin
    e0_G4_mul4_G16_inv0_G256_inv0_reg59 <= axorb_0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk60;
  assign clk60 = dec_255[0] & clk;

  always @(posedge clk60) begin
    e0_G4_mul4_G16_inv0_G256_inv0_reg60 <= cxord_0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk61;
  assign clk61 = ~dec_255[0] & clk;

  always @(posedge clk61) begin
    e0_G4_mul4_G16_inv0_G256_inv0_reg61 <= t309_axorb_0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk62;
  assign clk62 = ~dec_255[0] & clk;

  always @(posedge clk62) begin
    e0_G4_mul4_G16_inv0_G256_inv0_reg62 <= t326_cxord_0_G4_mul4_G16_inv0_G256_inv0;
  end

  assign t345_c0xord0_G16_inv0_G256_inv0 = y_reg247 ^ d0_G16_inv0_G256_inv0;
  assign t346_dec_1_inp = ~(~dec_1);
  assign t344_b0_G4_sq3_G16_inv0_G256_inv0 = ~(~t345_c0xord0_G16_inv0_G256_inv0 | y_reg249);
  assign t347_dec_1_inp = dec_1;
  assign t343_b0ls1_G4_sq3_G16_inv0_G256_inv0 = ~(~(t344_b0_G4_sq3_G16_inv0_G256_inv0 << y_reg251));
  assign t350_c0xord0_G16_inv0_G256_inv0 = y_reg252 ^ d0_G16_inv0_G256_inv0;
  assign t351_dec_2_inp = dec_2;
  assign t349_a0_0_G4_sq3_G16_inv0_G256_inv0 = ~(~t350_c0xord0_G16_inv0_G256_inv0 | y_reg254);
  assign t352_dec_1_inp = ~(~dec_1);
  assign t348_a0_G4_sq3_G16_inv0_G256_inv0 = ~(~(t349_a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg256));
  assign t342_e0_G16_inv0_G256_inv0 = ~(~t343_b0ls1_G4_sq3_G16_inv0_G256_inv0 & ~t348_a0_G4_sq3_G16_inv0_G256_inv0);
  assign t353_dec_1_inp = dec_1;
  assign t341_b0_G4_mul4_G16_inv0_G256_inv0 = ~t342_e0_G16_inv0_G256_inv0 | y_reg258;
  assign t358_p0ls2_G16_sq_scl0_G256_inv0 = p0_G16_sq_scl0_G256_inv0 << dec_2_inp;
  assign t359_q0_G16_sq_scl0_G256_inv0 = p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
  assign t357_c0_G256_inv0 = t358_p0ls2_G16_sq_scl0_G256_inv0 | t359_q0_G16_sq_scl0_G256_inv0;
  assign t361_p0ls2_G16_mul0_G256_inv0 = ~(~(p0_G16_mul0_G256_inv0 << y_reg259));
  assign t362_q0_G16_mul0_G256_inv0 = ~(~q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
  assign t360_d0_G256_inv0 = ~(~t361_p0ls2_G16_mul0_G256_inv0 & ~t362_q0_G16_mul0_G256_inv0);
  assign t356_c0xord0_G256_inv0 = ~(y_reg260 ^ ~t360_d0_G256_inv0);
  assign t363_dec_3_inp = dec_3;
  assign t355_b0_G16_inv0_G256_inv0 = ~(~t356_c0xord0_G256_inv0 | y_reg261);
  assign t364_dec_1_inp = dec_1;
  assign t354_d0_G4_mul4_G16_inv0_G256_inv0 = ~t355_b0_G16_inv0_G256_inv0 | y_reg262;
  wire clk63;
  assign clk63 = dec_45[1] & clk;

  always @(posedge clk63) begin
    q0_0_G4_mul4_G16_inv0_G256_inv0_reg63 <= b0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk64;
  assign clk64 = dec_45[1] & clk;

  always @(posedge clk64) begin
    q0_0_G4_mul4_G16_inv0_G256_inv0_reg64 <= d0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk65;
  assign clk65 = ~dec_45[1] & clk;

  always @(posedge clk65) begin
    q0_0_G4_mul4_G16_inv0_G256_inv0_reg65 <= t341_b0_G4_mul4_G16_inv0_G256_inv0;
  end

  wire clk66;
  assign clk66 = ~dec_45[1] & clk;

  always @(posedge clk66) begin
    q0_0_G4_mul4_G16_inv0_G256_inv0_reg66 <= t354_d0_G4_mul4_G16_inv0_G256_inv0;
  end

  assign t369_b0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg269;
  assign t370_dec_1_inp = ~(~dec_1);
  assign t368_b0ls1_G4_sq3_G16_inv0_G256_inv0 = t369_b0_G4_sq3_G16_inv0_G256_inv0 << y_reg271;
  assign t372_a0_0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg273;
  assign t373_dec_1_inp = dec_1;
  assign t371_a0_G4_sq3_G16_inv0_G256_inv0 = t372_a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg275;
  assign t367_e0_G16_inv0_G256_inv0 = t368_b0ls1_G4_sq3_G16_inv0_G256_inv0 | t371_a0_G4_sq3_G16_inv0_G256_inv0;
  assign t374_dec_2_inp = ~(~dec_2);
  assign t366_a0_0_G4_mul5_G16_inv0_G256_inv0 = ~(~t367_e0_G16_inv0_G256_inv0 | y_reg277);
  assign t375_dec_1_inp = ~(~dec_1);
  assign t365_a0_G4_mul5_G16_inv0_G256_inv0 = ~(t366_a0_0_G4_mul5_G16_inv0_G256_inv0 >> y_reg279);
  assign t380_c0xord0_G256_inv0 = y_reg280 ^ d0_G256_inv0;
  assign t381_dec_12_inp = ~(~dec_12);
  assign t379_a0_0_G16_inv0_G256_inv0 = t380_c0xord0_G256_inv0 & y_reg281;
  assign t382_dec_2_inp = ~(~dec_2);
  assign t378_a0_G16_inv0_G256_inv0 = t379_a0_0_G16_inv0_G256_inv0 >> y_reg282;
  assign t383_dec_2_inp = dec_2;
  assign t377_c0_0_G4_mul5_G16_inv0_G256_inv0 = ~(~t378_a0_G16_inv0_G256_inv0 | y_reg283);
  assign t384_dec_1_inp = ~(~dec_1);
  assign t376_c0_G4_mul5_G16_inv0_G256_inv0 = ~(t377_c0_0_G4_mul5_G16_inv0_G256_inv0 >> y_reg284);
  wire clk67;
  assign clk67 = dec_99[0] & clk;

  always @(posedge clk67) begin
    p0_0_G4_mul5_G16_inv0_G256_inv0_reg67 <= a0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk68;
  assign clk68 = dec_99[0] & clk;

  always @(posedge clk68) begin
    p0_0_G4_mul5_G16_inv0_G256_inv0_reg68 <= c0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk69;
  assign clk69 = ~dec_99[0] & clk;

  always @(posedge clk69) begin
    p0_0_G4_mul5_G16_inv0_G256_inv0_reg69 <= t365_a0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk70;
  assign clk70 = ~dec_99[0] & clk;

  always @(posedge clk70) begin
    p0_0_G4_mul5_G16_inv0_G256_inv0_reg70 <= t376_c0_G4_mul5_G16_inv0_G256_inv0;
  end

  assign t389_b0ls1_G4_sq3_G16_inv0_G256_inv0 = ~(~(b0_G4_sq3_G16_inv0_G256_inv0 << y_reg294));
  assign t390_a0_G4_sq3_G16_inv0_G256_inv0 = ~(~(a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg296));
  assign t388_e0_G16_inv0_G256_inv0 = t389_b0ls1_G4_sq3_G16_inv0_G256_inv0 | t390_a0_G4_sq3_G16_inv0_G256_inv0;
  assign t391_dec_2_inp = ~(~dec_2);
  assign t387_a0_0_G4_mul5_G16_inv0_G256_inv0 = t388_e0_G16_inv0_G256_inv0 & y_reg298;
  assign t392_dec_1_inp = ~(~dec_1);
  assign t386_a0_G4_mul5_G16_inv0_G256_inv0 = ~(~(t387_a0_0_G4_mul5_G16_inv0_G256_inv0 >> y_reg300));
  assign t396_b0_G4_sq3_G16_inv0_G256_inv0 = ~(~c0xord0_G16_inv0_G256_inv0 | y_reg302);
  assign t397_dec_1_inp = ~(~dec_1);
  assign t395_b0ls1_G4_sq3_G16_inv0_G256_inv0 = t396_b0_G4_sq3_G16_inv0_G256_inv0 << y_reg304;
  assign t399_a0_0_G4_sq3_G16_inv0_G256_inv0 = c0xord0_G16_inv0_G256_inv0 & y_reg306;
  assign t400_dec_1_inp = dec_1;
  assign t398_a0_G4_sq3_G16_inv0_G256_inv0 = ~(~(t399_a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg308));
  assign t394_e0_G16_inv0_G256_inv0 = ~(~t395_b0ls1_G4_sq3_G16_inv0_G256_inv0 & ~t398_a0_G4_sq3_G16_inv0_G256_inv0);
  assign t401_dec_1_inp = dec_1;
  assign t393_b0_G4_mul5_G16_inv0_G256_inv0 = ~(~t394_e0_G16_inv0_G256_inv0 | y_reg310);
  assign t385_axorb_0_G4_mul5_G16_inv0_G256_inv0 = ~(~(~t386_a0_G4_mul5_G16_inv0_G256_inv0)) ^ t393_b0_G4_mul5_G16_inv0_G256_inv0;
  assign t406_a0_0_G16_inv0_G256_inv0 = c0xord0_G256_inv0 & y_reg311;
  assign t407_dec_2_inp = ~(~dec_2);
  assign t405_a0_G16_inv0_G256_inv0 = ~(~(t406_a0_0_G16_inv0_G256_inv0 >> y_reg312));
  assign t408_dec_2_inp = dec_2;
  assign t404_c0_0_G4_mul5_G16_inv0_G256_inv0 = t405_a0_G16_inv0_G256_inv0 & y_reg313;
  assign t409_dec_1_inp = dec_1;
  assign t403_c0_G4_mul5_G16_inv0_G256_inv0 = ~(~(t404_c0_0_G4_mul5_G16_inv0_G256_inv0 >> y_reg314));
  assign t413_c0xord0_G256_inv0 = ~(y_reg315 ^ d0_G256_inv0);
  assign t414_dec_12_inp = ~(~dec_12);
  assign t412_a0_0_G16_inv0_G256_inv0 = t413_c0xord0_G256_inv0 & y_reg316;
  assign t415_dec_2_inp = dec_2;
  assign t411_a0_G16_inv0_G256_inv0 = t412_a0_0_G16_inv0_G256_inv0 >> y_reg317;
  assign t416_dec_1_inp = dec_1;
  assign t410_d0_G4_mul5_G16_inv0_G256_inv0 = t411_a0_G16_inv0_G256_inv0 & y_reg318;
  assign t402_cxord_0_G4_mul5_G16_inv0_G256_inv0 = ~t403_c0_G4_mul5_G16_inv0_G256_inv0 ^ t410_d0_G4_mul5_G16_inv0_G256_inv0;
  wire clk71;
  assign clk71 = dec_3[1] & clk;

  always @(posedge clk71) begin
    e0_G4_mul5_G16_inv0_G256_inv0_reg71 <= a0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk72;
  assign clk72 = dec_3[1] & clk;

  always @(posedge clk72) begin
    e0_G4_mul5_G16_inv0_G256_inv0_reg72 <= b0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk73;
  assign clk73 = dec_3[1] & clk;

  always @(posedge clk73) begin
    e0_G4_mul5_G16_inv0_G256_inv0_reg73 <= c0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk74;
  assign clk74 = dec_3[1] & clk;

  always @(posedge clk74) begin
    e0_G4_mul5_G16_inv0_G256_inv0_reg74 <= d0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk75;
  assign clk75 = ~dec_3[1] & clk;

  always @(posedge clk75) begin
    e0_G4_mul5_G16_inv0_G256_inv0_reg75 <= t385_axorb_0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk76;
  assign clk76 = ~dec_3[1] & clk;

  always @(posedge clk76) begin
    e0_G4_mul5_G16_inv0_G256_inv0_reg76 <= t402_cxord_0_G4_mul5_G16_inv0_G256_inv0;
  end

  assign t421_c0xord0_G16_inv0_G256_inv0 = y_reg327 ^ d0_G16_inv0_G256_inv0;
  assign t422_dec_1_inp = ~(~dec_1);
  assign t420_b0_G4_sq3_G16_inv0_G256_inv0 = ~(~t421_c0xord0_G16_inv0_G256_inv0 | y_reg329);
  assign t423_dec_1_inp = dec_1;
  assign t419_b0ls1_G4_sq3_G16_inv0_G256_inv0 = t420_b0_G4_sq3_G16_inv0_G256_inv0 << y_reg331;
  assign t426_c0xord0_G16_inv0_G256_inv0 = y_reg332 ^ d0_G16_inv0_G256_inv0;
  assign t427_dec_2_inp = dec_2;
  assign t425_a0_0_G4_sq3_G16_inv0_G256_inv0 = ~(~t426_c0xord0_G16_inv0_G256_inv0 | y_reg334);
  assign t428_dec_1_inp = ~(~dec_1);
  assign t424_a0_G4_sq3_G16_inv0_G256_inv0 = t425_a0_0_G4_sq3_G16_inv0_G256_inv0 >> y_reg336;
  assign t418_e0_G16_inv0_G256_inv0 = ~t419_b0ls1_G4_sq3_G16_inv0_G256_inv0 & ~t424_a0_G4_sq3_G16_inv0_G256_inv0;
  assign t429_dec_1_inp = ~dec_1;
  assign t417_b0_G4_mul5_G16_inv0_G256_inv0 = t418_e0_G16_inv0_G256_inv0 | y_reg338;
  assign t434_c0_G256_inv0 = p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0;
  assign t435_d0_G256_inv0 = ~(~p0ls2_G16_mul0_G256_inv0 & ~q0_G16_mul0_G256_inv0);
  assign t433_c0xord0_G256_inv0 = ~(y_reg339 ^ ~t435_d0_G256_inv0);
  assign t436_dec_12_inp = dec_12;
  assign t432_a0_0_G16_inv0_G256_inv0 = ~(~t433_c0xord0_G256_inv0 | y_reg340);
  assign t437_dec_2_inp = dec_2;
  assign t431_a0_G16_inv0_G256_inv0 = ~(t432_a0_0_G16_inv0_G256_inv0 >> y_reg341);
  assign t438_dec_1_inp = ~dec_1;
  assign t430_d0_G4_mul5_G16_inv0_G256_inv0 = t431_a0_G16_inv0_G256_inv0 | y_reg342;
  wire clk77;
  assign clk77 = dec_9[1] & clk;

  always @(posedge clk77) begin
    q0_0_G4_mul5_G16_inv0_G256_inv0_reg77 <= b0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk78;
  assign clk78 = dec_9[1] & clk;

  always @(posedge clk78) begin
    q0_0_G4_mul5_G16_inv0_G256_inv0_reg78 <= d0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk79;
  assign clk79 = ~dec_9[1] & clk;

  always @(posedge clk79) begin
    q0_0_G4_mul5_G16_inv0_G256_inv0_reg79 <= t417_b0_G4_mul5_G16_inv0_G256_inv0;
  end

  wire clk80;
  assign clk80 = ~dec_9[1] & clk;

  always @(posedge clk80) begin
    q0_0_G4_mul5_G16_inv0_G256_inv0_reg80 <= t430_d0_G4_mul5_G16_inv0_G256_inv0;
  end

  assign t443_a0_0_G16_mul1_G256_inv0 = ~(~e0_G256_inv0 | y_reg429);
  assign t444_dec_2_inp = dec_2;
  assign t442_a0_G16_mul1_G256_inv0 = ~(~(t443_a0_0_G16_mul1_G256_inv0 >> y_reg432));
  assign t446_e0_G256_inv0 = ~(~p0ls2_G16_inv0_G256_inv0 & ~q0_G16_inv0_G256_inv0);
  assign t447_dec_3_inp = dec_3;
  assign t445_b0_G16_mul1_G256_inv0 = t446_e0_G256_inv0 & y_reg435;
  assign t441_axorb_0_G16_mul1_G256_inv0 = ~(~t442_a0_G16_mul1_G256_inv0 ^ t445_b0_G16_mul1_G256_inv0);
  assign t448_dec_2_inp = ~(~dec_2);
  assign t440_a0_0_G4_mul0_G16_mul1_G256_inv0 = ~(~t441_axorb_0_G16_mul1_G256_inv0 | y_reg438);
  assign t449_dec_1_inp = dec_1;
  assign t439_a0_G4_mul0_G16_mul1_G256_inv0 = ~(t440_a0_0_G4_mul0_G16_mul1_G256_inv0 >> y_reg441);
  assign t454_c0_0_G16_mul1_G256_inv0 = b0_G256_inv0 & dec_12_inp;
  assign t455_dec_2_inp = ~(~dec_2);
  assign t453_c0_G16_mul1_G256_inv0 = t454_c0_0_G16_mul1_G256_inv0 >> t455_dec_2_inp;
  assign t457_b0_G256_inv0 = ~(~t2 | ~dec_15_inp);
  assign t458_dec_3_inp = dec_3;
  assign t456_d0_G16_mul1_G256_inv0 = ~(~t457_b0_G256_inv0 | ~t458_dec_3_inp);
  assign t452_cxord_0_G16_mul1_G256_inv0 = ~(~t453_c0_G16_mul1_G256_inv0 ^ t456_d0_G16_mul1_G256_inv0);
  assign t459_dec_2_inp = dec_2;
  assign t451_c0_0_G4_mul0_G16_mul1_G256_inv0 = t452_cxord_0_G16_mul1_G256_inv0 & t459_dec_2_inp;
  assign t460_dec_1_inp = dec_1;
  assign t450_c0_G4_mul0_G16_mul1_G256_inv0 = ~(t451_c0_0_G4_mul0_G16_mul1_G256_inv0 >> t460_dec_1_inp);
  wire clk81;
  assign clk81 = dec_11[2] & clk;

  always @(posedge clk81) begin
    p0_0_G4_mul0_G16_mul1_G256_inv0_reg81 <= a0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk82;
  assign clk82 = dec_11[2] & clk;

  always @(posedge clk82) begin
    p0_0_G4_mul0_G16_mul1_G256_inv0_reg82 <= c0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk83;
  assign clk83 = ~dec_11[2] & clk;

  always @(posedge clk83) begin
    p0_0_G4_mul0_G16_mul1_G256_inv0_reg83 <= t439_a0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk84;
  assign clk84 = ~dec_11[2] & clk;

  always @(posedge clk84) begin
    p0_0_G4_mul0_G16_mul1_G256_inv0_reg84 <= t450_c0_G4_mul0_G16_mul1_G256_inv0;
  end

  assign t465_a0_G16_mul1_G256_inv0 = a0_0_G16_mul1_G256_inv0 >> y_reg459;
  assign t466_b0_G16_mul1_G256_inv0 = e0_G256_inv0 & y_reg462;
  assign t464_axorb_0_G16_mul1_G256_inv0 = t465_a0_G16_mul1_G256_inv0 ^ t466_b0_G16_mul1_G256_inv0;
  assign t467_dec_2_inp = ~(~dec_2);
  assign t463_a0_0_G4_mul0_G16_mul1_G256_inv0 = t464_axorb_0_G16_mul1_G256_inv0 & y_reg465;
  assign t468_dec_1_inp = ~(~dec_1);
  assign t462_a0_G4_mul0_G16_mul1_G256_inv0 = ~(~(t463_a0_0_G4_mul0_G16_mul1_G256_inv0 >> y_reg468));
  assign t472_a0_0_G16_mul1_G256_inv0 = ~(~e0_G256_inv0 | y_reg471);
  assign t473_dec_2_inp = ~(~dec_2);
  assign t471_a0_G16_mul1_G256_inv0 = t472_a0_0_G16_mul1_G256_inv0 >> y_reg474;
  assign t475_e0_G256_inv0 = ~(~p0ls2_G16_inv0_G256_inv0 & ~q0_G16_inv0_G256_inv0);
  assign t476_dec_3_inp = ~(~dec_3);
  assign t474_b0_G16_mul1_G256_inv0 = t475_e0_G256_inv0 & y_reg477;
  assign t470_axorb_0_G16_mul1_G256_inv0 = t471_a0_G16_mul1_G256_inv0 ^ t474_b0_G16_mul1_G256_inv0;
  assign t477_dec_1_inp = dec_1;
  assign t469_b0_G4_mul0_G16_mul1_G256_inv0 = ~(~t470_axorb_0_G16_mul1_G256_inv0 | y_reg480);
  assign t461_axorb_0_G4_mul0_G16_mul1_G256_inv0 = ~(~t462_a0_G4_mul0_G16_mul1_G256_inv0) ^ ~t469_b0_G4_mul0_G16_mul1_G256_inv0;
  assign t482_c0_G16_mul1_G256_inv0 = c0_0_G16_mul1_G256_inv0 >> dec_2_inp;
  assign t483_d0_G16_mul1_G256_inv0 = ~(~b0_G256_inv0 | ~dec_3_inp);
  assign t481_cxord_0_G16_mul1_G256_inv0 = ~(t482_c0_G16_mul1_G256_inv0 ^ ~t483_d0_G16_mul1_G256_inv0);
  assign t484_dec_2_inp = dec_2;
  assign t480_c0_0_G4_mul0_G16_mul1_G256_inv0 = ~(~t481_cxord_0_G16_mul1_G256_inv0 | ~t484_dec_2_inp);
  assign t485_dec_1_inp = ~(~dec_1);
  assign t479_c0_G4_mul0_G16_mul1_G256_inv0 = t480_c0_0_G4_mul0_G16_mul1_G256_inv0 >> t485_dec_1_inp;
  assign t489_c0_0_G16_mul1_G256_inv0 = b0_G256_inv0 & dec_12_inp;
  assign t490_dec_2_inp = ~(~dec_2);
  assign t488_c0_G16_mul1_G256_inv0 = ~(~(t489_c0_0_G16_mul1_G256_inv0 >> t490_dec_2_inp));
  assign t492_b0_G256_inv0 = t2 & dec_15_inp;
  assign t493_dec_3_inp = ~(~dec_3);
  assign t491_d0_G16_mul1_G256_inv0 = t492_b0_G256_inv0 & t493_dec_3_inp;
  assign t487_cxord_0_G16_mul1_G256_inv0 = ~(t488_c0_G16_mul1_G256_inv0 ^ ~t491_d0_G16_mul1_G256_inv0);
  assign t494_dec_1_inp = dec_1;
  assign t486_d0_G4_mul0_G16_mul1_G256_inv0 = t487_cxord_0_G16_mul1_G256_inv0 & t494_dec_1_inp;
  assign t478_cxord_0_G4_mul0_G16_mul1_G256_inv0 = ~t479_c0_G4_mul0_G16_mul1_G256_inv0 ^ t486_d0_G4_mul0_G16_mul1_G256_inv0;
  wire clk85;
  assign clk85 = dec_36[7] & clk;

  always @(posedge clk85) begin
    e0_G4_mul0_G16_mul1_G256_inv0_reg85 <= a0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk86;
  assign clk86 = dec_36[7] & clk;

  always @(posedge clk86) begin
    e0_G4_mul0_G16_mul1_G256_inv0_reg86 <= b0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk87;
  assign clk87 = dec_36[7] & clk;

  always @(posedge clk87) begin
    e0_G4_mul0_G16_mul1_G256_inv0_reg87 <= c0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk88;
  assign clk88 = dec_36[7] & clk;

  always @(posedge clk88) begin
    e0_G4_mul0_G16_mul1_G256_inv0_reg88 <= d0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk89;
  assign clk89 = ~dec_36[7] & clk;

  always @(posedge clk89) begin
    e0_G4_mul0_G16_mul1_G256_inv0_reg89 <= t461_axorb_0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk90;
  assign clk90 = ~dec_36[7] & clk;

  always @(posedge clk90) begin
    e0_G4_mul0_G16_mul1_G256_inv0_reg90 <= t478_cxord_0_G4_mul0_G16_mul1_G256_inv0;
  end

  assign t499_e0_G256_inv0 = p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0;
  assign t500_dec_12_inp = ~(~dec_12);
  assign t498_a0_0_G16_mul1_G256_inv0 = t499_e0_G256_inv0 & y_reg496;
  assign t501_dec_2_inp = dec_2;
  assign t497_a0_G16_mul1_G256_inv0 = t498_a0_0_G16_mul1_G256_inv0 >> y_reg499;
  assign t504_p0ls2_G16_inv0_G256_inv0 = ~(~(p0_G16_inv0_G256_inv0 << y_reg502));
  assign t505_q0_G16_inv0_G256_inv0 = p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0;
  assign t503_e0_G256_inv0 = ~(~t504_p0ls2_G16_inv0_G256_inv0 & ~t505_q0_G16_inv0_G256_inv0);
  assign t506_dec_3_inp = dec_3;
  assign t502_b0_G16_mul1_G256_inv0 = ~(~t503_e0_G256_inv0 | y_reg505);
  assign t496_axorb_0_G16_mul1_G256_inv0 = ~(t497_a0_G16_mul1_G256_inv0 ^ ~t502_b0_G16_mul1_G256_inv0);
  assign t507_dec_1_inp = ~(~dec_1);
  assign t495_b0_G4_mul0_G16_mul1_G256_inv0 = t496_axorb_0_G16_mul1_G256_inv0 & y_reg508;
  assign t512_b0_G256_inv0 = ~(~t2 | ~dec_15_inp);
  assign t513_dec_12_inp = ~(~dec_12);
  assign t511_c0_0_G16_mul1_G256_inv0 = t512_b0_G256_inv0 & t513_dec_12_inp;
  assign t514_dec_2_inp = dec_2;
  assign t510_c0_G16_mul1_G256_inv0 = t511_c0_0_G16_mul1_G256_inv0 >> t514_dec_2_inp;
  assign t518_y8_G256_newbasis0 = ~(~ny8_G256_newbasis0 + (~tempyIntoNegCond8_G256_newbasis0 + 1));
  assign t517_t2 = ~(~t518_y8_G256_newbasis0);
  assign t519_dec_15_inp = dec_15;
  assign t516_b0_G256_inv0 = t517_t2 & t519_dec_15_inp;
  assign t520_dec_3_inp = ~(~dec_3);
  assign t515_d0_G16_mul1_G256_inv0 = t516_b0_G256_inv0 & t520_dec_3_inp;
  assign t509_cxord_0_G16_mul1_G256_inv0 = t510_c0_G16_mul1_G256_inv0 ^ t515_d0_G16_mul1_G256_inv0;
  assign t521_dec_1_inp = ~(~dec_1);
  assign t508_d0_G4_mul0_G16_mul1_G256_inv0 = ~(~t509_cxord_0_G16_mul1_G256_inv0 | ~t521_dec_1_inp);
  wire clk91;
  assign clk91 = dec_12[3] & clk;

  always @(posedge clk91) begin
    q0_0_G4_mul0_G16_mul1_G256_inv0_reg91 <= b0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk92;
  assign clk92 = dec_12[3] & clk;

  always @(posedge clk92) begin
    q0_0_G4_mul0_G16_mul1_G256_inv0_reg92 <= d0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk93;
  assign clk93 = ~dec_12[3] & clk;

  always @(posedge clk93) begin
    q0_0_G4_mul0_G16_mul1_G256_inv0_reg93 <= t495_b0_G4_mul0_G16_mul1_G256_inv0;
  end

  wire clk94;
  assign clk94 = ~dec_12[3] & clk;

  always @(posedge clk94) begin
    q0_0_G4_mul0_G16_mul1_G256_inv0_reg94 <= t508_d0_G4_mul0_G16_mul1_G256_inv0;
  end

  assign t526_e0_G256_inv0 = ~(~p0ls2_G16_inv0_G256_inv0 & ~q0_G16_inv0_G256_inv0);
  assign t527_dec_12_inp = dec_12;
  assign t525_a0_0_G16_mul1_G256_inv0 = t526_e0_G256_inv0 & y_reg347;
  assign t528_dec_2_inp = ~(~dec_2);
  assign t524_a0_G16_mul1_G256_inv0 = ~(~(t525_a0_0_G16_mul1_G256_inv0 >> y_reg350));
  assign t529_dec_2_inp = ~(~dec_2);
  assign t523_a0_0_G4_mul1_G16_mul1_G256_inv0 = t524_a0_G16_mul1_G256_inv0 & y_reg353;
  assign t530_dec_1_inp = ~(~dec_1);
  assign t522_a0_G4_mul1_G16_mul1_G256_inv0 = ~(t523_a0_0_G4_mul1_G16_mul1_G256_inv0 >> y_reg356);
  assign t535_b0_G256_inv0 = t2 & dec_15_inp;
  assign t536_dec_12_inp = ~(~dec_12);
  assign t534_c0_0_G16_mul1_G256_inv0 = ~(~t535_b0_G256_inv0 | ~t536_dec_12_inp);
  assign t537_dec_2_inp = dec_2;
  assign t533_c0_G16_mul1_G256_inv0 = t534_c0_0_G16_mul1_G256_inv0 >> t537_dec_2_inp;
  assign t538_dec_2_inp = dec_2;
  assign t532_c0_0_G4_mul1_G16_mul1_G256_inv0 = t533_c0_G16_mul1_G256_inv0 & t538_dec_2_inp;
  assign t539_dec_1_inp = ~(~dec_1);
  assign t531_c0_G4_mul1_G16_mul1_G256_inv0 = ~(t532_c0_0_G4_mul1_G16_mul1_G256_inv0 >> t539_dec_1_inp);
  wire clk95;
  assign clk95 = dec_1[1] & clk;

  always @(posedge clk95) begin
    p0_0_G4_mul1_G16_mul1_G256_inv0_reg95 <= a0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk96;
  assign clk96 = dec_1[1] & clk;

  always @(posedge clk96) begin
    p0_0_G4_mul1_G16_mul1_G256_inv0_reg96 <= c0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk97;
  assign clk97 = ~dec_1[1] & clk;

  always @(posedge clk97) begin
    p0_0_G4_mul1_G16_mul1_G256_inv0_reg97 <= t522_a0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk98;
  assign clk98 = ~dec_1[1] & clk;

  always @(posedge clk98) begin
    p0_0_G4_mul1_G16_mul1_G256_inv0_reg98 <= t531_c0_G4_mul1_G16_mul1_G256_inv0;
  end

  assign t544_a0_0_G16_mul1_G256_inv0 = ~(~e0_G256_inv0 | y_reg377);
  assign t545_dec_2_inp = dec_2;
  assign t543_a0_G16_mul1_G256_inv0 = t544_a0_0_G16_mul1_G256_inv0 >> y_reg380;
  assign t546_dec_2_inp = dec_2;
  assign t542_a0_0_G4_mul1_G16_mul1_G256_inv0 = ~(~t543_a0_G16_mul1_G256_inv0 | y_reg383);
  assign t547_dec_1_inp = ~(~dec_1);
  assign t541_a0_G4_mul1_G16_mul1_G256_inv0 = ~(~(t542_a0_0_G4_mul1_G16_mul1_G256_inv0 >> y_reg386));
  assign t551_e0_G256_inv0 = p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0;
  assign t552_dec_12_inp = dec_12;
  assign t550_a0_0_G16_mul1_G256_inv0 = ~(~t551_e0_G256_inv0 | y_reg389);
  assign t553_dec_2_inp = dec_2;
  assign t549_a0_G16_mul1_G256_inv0 = t550_a0_0_G16_mul1_G256_inv0 >> y_reg392;
  assign t554_dec_1_inp = ~(~dec_1);
  assign t548_b0_G4_mul1_G16_mul1_G256_inv0 = ~(~t549_a0_G16_mul1_G256_inv0 | y_reg395);
  assign t540_axorb_0_G4_mul1_G16_mul1_G256_inv0 = ~t541_a0_G4_mul1_G16_mul1_G256_inv0 ^ t548_b0_G4_mul1_G16_mul1_G256_inv0;
  assign t559_c0_0_G16_mul1_G256_inv0 = b0_G256_inv0 & dec_12_inp;
  assign t560_dec_2_inp = dec_2;
  assign t558_c0_G16_mul1_G256_inv0 = ~(~(t559_c0_0_G16_mul1_G256_inv0 >> t560_dec_2_inp));
  assign t561_dec_2_inp = ~(~dec_2);
  assign t557_c0_0_G4_mul1_G16_mul1_G256_inv0 = t558_c0_G16_mul1_G256_inv0 & t561_dec_2_inp;
  assign t562_dec_1_inp = dec_1;
  assign t556_c0_G4_mul1_G16_mul1_G256_inv0 = ~(~(t557_c0_0_G4_mul1_G16_mul1_G256_inv0 >> t562_dec_1_inp));
  assign t566_b0_G256_inv0 = t2 & dec_15_inp;
  assign t567_dec_12_inp = ~(~dec_12);
  assign t565_c0_0_G16_mul1_G256_inv0 = t566_b0_G256_inv0 & t567_dec_12_inp;
  assign t568_dec_2_inp = dec_2;
  assign t564_c0_G16_mul1_G256_inv0 = ~(~(t565_c0_0_G16_mul1_G256_inv0 >> t568_dec_2_inp));
  assign t569_dec_1_inp = ~(~dec_1);
  assign t563_d0_G4_mul1_G16_mul1_G256_inv0 = ~(~t564_c0_G16_mul1_G256_inv0 | ~t569_dec_1_inp);
  assign t555_cxord_0_G4_mul1_G16_mul1_G256_inv0 = ~t556_c0_G4_mul1_G16_mul1_G256_inv0 ^ ~(~t563_d0_G4_mul1_G16_mul1_G256_inv0);
  wire clk99;
  assign clk99 = dec_88[0] & clk;

  always @(posedge clk99) begin
    e0_G4_mul1_G16_mul1_G256_inv0_reg99 <= a0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk100;
  assign clk100 = dec_88[0] & clk;

  always @(posedge clk100) begin
    e0_G4_mul1_G16_mul1_G256_inv0_reg100 <= b0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk101;
  assign clk101 = dec_88[0] & clk;

  always @(posedge clk101) begin
    e0_G4_mul1_G16_mul1_G256_inv0_reg101 <= c0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk102;
  assign clk102 = dec_88[0] & clk;

  always @(posedge clk102) begin
    e0_G4_mul1_G16_mul1_G256_inv0_reg102 <= d0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk103;
  assign clk103 = ~dec_88[0] & clk;

  always @(posedge clk103) begin
    e0_G4_mul1_G16_mul1_G256_inv0_reg103 <= t540_axorb_0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk104;
  assign clk104 = ~dec_88[0] & clk;

  always @(posedge clk104) begin
    e0_G4_mul1_G16_mul1_G256_inv0_reg104 <= t555_cxord_0_G4_mul1_G16_mul1_G256_inv0;
  end

  assign t574_p0ls2_G16_inv0_G256_inv0 = p0_G16_inv0_G256_inv0 << y_reg411;
  assign t575_q0_G16_inv0_G256_inv0 = p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0;
  assign t573_e0_G256_inv0 = ~(~t574_p0ls2_G16_inv0_G256_inv0 & ~t575_q0_G16_inv0_G256_inv0);
  assign t576_dec_12_inp = ~(~dec_12);
  assign t572_a0_0_G16_mul1_G256_inv0 = ~(~t573_e0_G256_inv0 | y_reg414);
  assign t577_dec_2_inp = dec_2;
  assign t571_a0_G16_mul1_G256_inv0 = ~(~(t572_a0_0_G16_mul1_G256_inv0 >> y_reg417));
  assign t578_dec_1_inp = dec_1;
  assign t570_b0_G4_mul1_G16_mul1_G256_inv0 = ~t571_a0_G16_mul1_G256_inv0 | y_reg420;
  assign t584_y8_G256_newbasis0 = ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0;
  assign t583_t2 = ~(~t584_y8_G256_newbasis0);
  assign t585_dec_15_inp = dec_15;
  assign t582_b0_G256_inv0 = t583_t2 & t585_dec_15_inp;
  assign t586_dec_12_inp = ~(~dec_12);
  assign t581_c0_0_G16_mul1_G256_inv0 = ~(~t582_b0_G256_inv0 | ~t586_dec_12_inp);
  assign t587_dec_2_inp = ~(~dec_2);
  assign t580_c0_G16_mul1_G256_inv0 = ~(t581_c0_0_G16_mul1_G256_inv0 >> t587_dec_2_inp);
  assign t588_dec_1_inp = ~dec_1;
  assign t579_d0_G4_mul1_G16_mul1_G256_inv0 = t580_c0_G16_mul1_G256_inv0 | t588_dec_1_inp;
  wire clk105;
  assign clk105 = dec_3[1] & clk;

  always @(posedge clk105) begin
    q0_0_G4_mul1_G16_mul1_G256_inv0_reg105 <= b0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk106;
  assign clk106 = dec_3[1] & clk;

  always @(posedge clk106) begin
    q0_0_G4_mul1_G16_mul1_G256_inv0_reg106 <= d0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk107;
  assign clk107 = ~dec_3[1] & clk;

  always @(posedge clk107) begin
    q0_0_G4_mul1_G16_mul1_G256_inv0_reg107 <= t570_b0_G4_mul1_G16_mul1_G256_inv0;
  end

  wire clk108;
  assign clk108 = ~dec_3[1] & clk;

  always @(posedge clk108) begin
    q0_0_G4_mul1_G16_mul1_G256_inv0_reg108 <= t579_d0_G4_mul1_G16_mul1_G256_inv0;
  end

  assign t593_p0ls2_G16_inv0_G256_inv0 = ~(~(p0_G16_inv0_G256_inv0 << y_reg537));
  assign t594_q0_G16_inv0_G256_inv0 = p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0;
  assign t592_e0_G256_inv0 = t593_p0ls2_G16_inv0_G256_inv0 | t594_q0_G16_inv0_G256_inv0;
  assign t595_dec_3_inp = dec_3;
  assign t591_b0_G16_mul1_G256_inv0 = ~(~t592_e0_G256_inv0 | y_reg540);
  assign t596_dec_2_inp = ~(~dec_2);
  assign t590_a0_0_G4_mul2_G16_mul1_G256_inv0 = ~(~t591_b0_G16_mul1_G256_inv0 | y_reg543);
  assign t597_dec_1_inp = ~(~dec_1);
  assign t589_a0_G4_mul2_G16_mul1_G256_inv0 = ~(t590_a0_0_G4_mul2_G16_mul1_G256_inv0 >> y_reg546);
  assign t603_y8_G256_newbasis0 = ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0;
  assign t602_t2 = ~(~t603_y8_G256_newbasis0);
  assign t604_dec_15_inp = dec_15;
  assign t601_b0_G256_inv0 = ~(~t602_t2 | ~t604_dec_15_inp);
  assign t605_dec_3_inp = dec_3;
  assign t600_d0_G16_mul1_G256_inv0 = ~(~t601_b0_G256_inv0 | ~t605_dec_3_inp);
  assign t606_dec_2_inp = dec_2;
  assign t599_c0_0_G4_mul2_G16_mul1_G256_inv0 = ~(~t600_d0_G16_mul1_G256_inv0 | ~t606_dec_2_inp);
  assign t607_dec_1_inp = dec_1;
  assign t598_c0_G4_mul2_G16_mul1_G256_inv0 = ~(t599_c0_0_G4_mul2_G16_mul1_G256_inv0 >> t607_dec_1_inp);
  wire clk109;
  assign clk109 = r[19] & clk;

  always @(posedge clk109) begin
    p0_0_G4_mul2_G16_mul1_G256_inv0_reg109 <= a0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk110;
  assign clk110 = r[19] & clk;

  always @(posedge clk110) begin
    p0_0_G4_mul2_G16_mul1_G256_inv0_reg110 <= c0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk111;
  assign clk111 = ~r[19] & clk;

  always @(posedge clk111) begin
    p0_0_G4_mul2_G16_mul1_G256_inv0_reg111 <= t589_a0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk112;
  assign clk112 = ~r[19] & clk;

  always @(posedge clk112) begin
    p0_0_G4_mul2_G16_mul1_G256_inv0_reg112 <= t598_c0_G4_mul2_G16_mul1_G256_inv0;
  end

  assign t612_e0_G256_inv0 = p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0;
  assign t613_dec_3_inp = ~(~dec_3);
  assign t611_b0_G16_mul1_G256_inv0 = t612_e0_G256_inv0 & y_reg561;
  assign t614_dec_2_inp = dec_2;
  assign t610_a0_0_G4_mul2_G16_mul1_G256_inv0 = ~(~t611_b0_G16_mul1_G256_inv0 | y_reg564);
  assign t615_dec_1_inp = dec_1;
  assign t609_a0_G4_mul2_G16_mul1_G256_inv0 = ~(~(t610_a0_0_G4_mul2_G16_mul1_G256_inv0 >> y_reg567));
  assign t619_p0ls2_G16_inv0_G256_inv0 = ~(~(p0_G16_inv0_G256_inv0 << y_reg570));
  assign t620_q0_G16_inv0_G256_inv0 = ~(~p0ls1_G4_mul5_G16_inv0_G256_inv0 & ~q0_G4_mul5_G16_inv0_G256_inv0);
  assign t618_e0_G256_inv0 = t619_p0ls2_G16_inv0_G256_inv0 | t620_q0_G16_inv0_G256_inv0;
  assign t621_dec_3_inp = dec_3;
  assign t617_b0_G16_mul1_G256_inv0 = ~(~t618_e0_G256_inv0 | y_reg573);
  assign t622_dec_1_inp = ~(~dec_1);
  assign t616_b0_G4_mul2_G16_mul1_G256_inv0 = ~t617_b0_G16_mul1_G256_inv0 | y_reg576;
  assign t608_axorb_0_G4_mul2_G16_mul1_G256_inv0 = ~t609_a0_G4_mul2_G16_mul1_G256_inv0 ^ ~t616_b0_G4_mul2_G16_mul1_G256_inv0;
  assign t627_b0_G256_inv0 = t2 & dec_15_inp;
  assign t628_dec_3_inp = dec_3;
  assign t626_d0_G16_mul1_G256_inv0 = t627_b0_G256_inv0 & t628_dec_3_inp;
  assign t629_dec_2_inp = dec_2;
  assign t625_c0_0_G4_mul2_G16_mul1_G256_inv0 = t626_d0_G16_mul1_G256_inv0 & t629_dec_2_inp;
  assign t630_dec_1_inp = ~(~dec_1);
  assign t624_c0_G4_mul2_G16_mul1_G256_inv0 = ~(~(t625_c0_0_G4_mul2_G16_mul1_G256_inv0 >> t630_dec_1_inp));
  assign t635_y8_G256_newbasis0 = ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0;
  assign t634_t2 = t635_y8_G256_newbasis0;
  assign t636_dec_15_inp = ~(~dec_15);
  assign t633_b0_G256_inv0 = ~(~t634_t2 | ~t636_dec_15_inp);
  assign t637_dec_3_inp = dec_3;
  assign t632_d0_G16_mul1_G256_inv0 = ~t633_b0_G256_inv0 | ~t637_dec_3_inp;
  assign t638_dec_1_inp = ~dec_1;
  assign t631_d0_G4_mul2_G16_mul1_G256_inv0 = t632_d0_G16_mul1_G256_inv0 | t638_dec_1_inp;
  assign t623_cxord_0_G4_mul2_G16_mul1_G256_inv0 = ~t624_c0_G4_mul2_G16_mul1_G256_inv0 ^ ~t631_d0_G4_mul2_G16_mul1_G256_inv0;
  wire clk113;
  assign clk113 = dec_11[2] & clk;

  always @(posedge clk113) begin
    e0_G4_mul2_G16_mul1_G256_inv0_reg113 <= axorb_0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk114;
  assign clk114 = dec_11[2] & clk;

  always @(posedge clk114) begin
    e0_G4_mul2_G16_mul1_G256_inv0_reg114 <= cxord_0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk115;
  assign clk115 = ~dec_11[2] & clk;

  always @(posedge clk115) begin
    e0_G4_mul2_G16_mul1_G256_inv0_reg115 <= t608_axorb_0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk116;
  assign clk116 = ~dec_11[2] & clk;

  always @(posedge clk116) begin
    e0_G4_mul2_G16_mul1_G256_inv0_reg116 <= t623_cxord_0_G4_mul2_G16_mul1_G256_inv0;
  end

  assign t643_p0_G16_inv0_G256_inv0 = ~(~p0ls1_G4_mul4_G16_inv0_G256_inv0 & ~q0_G4_mul4_G16_inv0_G256_inv0);
  assign t644_dec_2_inp = ~(~dec_2);
  assign t642_p0ls2_G16_inv0_G256_inv0 = t643_p0_G16_inv0_G256_inv0 << y_reg592;
  assign t646_p0ls1_G4_mul5_G16_inv0_G256_inv0 = ~(~(p0_G4_mul5_G16_inv0_G256_inv0 << y_reg595));
  assign t647_q0_G4_mul5_G16_inv0_G256_inv0 = q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0;
  assign t645_q0_G16_inv0_G256_inv0 = ~(~t646_p0ls1_G4_mul5_G16_inv0_G256_inv0 & ~t647_q0_G4_mul5_G16_inv0_G256_inv0);
  assign t641_e0_G256_inv0 = ~(~t642_p0ls2_G16_inv0_G256_inv0 & ~t645_q0_G16_inv0_G256_inv0);
  assign t648_dec_3_inp = dec_3;
  assign t640_b0_G16_mul1_G256_inv0 = t641_e0_G256_inv0 & y_reg598;
  assign t649_dec_1_inp = dec_1;
  assign t639_b0_G4_mul2_G16_mul1_G256_inv0 = ~t640_b0_G16_mul1_G256_inv0 | y_reg601;
  assign t655_ny8_G256_newbasis0 = cond8_G256_newbasis0 * yxorb8_G256_newbasis0;
  assign t656_tempyIntoNegCond8_G256_newbasis0 = ~((~(tempy8_G256_newbasis0 + negCond8_G256_newbasis0) << 7 + 1) - ~tempy8_G256_newbasis0 * ~negCond8_G256_newbasis0 + (tempy8_G256_newbasis0 + negCond8_G256_newbasis0));
  assign t654_y8_G256_newbasis0 = ~(~t655_ny8_G256_newbasis0 + (~t656_tempyIntoNegCond8_G256_newbasis0 + 1));
  assign t653_t2 = t654_y8_G256_newbasis0;
  assign t657_dec_15_inp = dec_15;
  assign t652_b0_G256_inv0 = ~(~t653_t2 | ~t657_dec_15_inp);
  assign t658_dec_3_inp = dec_3;
  assign t651_d0_G16_mul1_G256_inv0 = ~(~t652_b0_G256_inv0 | ~t658_dec_3_inp);
  assign t659_dec_1_inp = dec_1;
  assign t650_d0_G4_mul2_G16_mul1_G256_inv0 = ~t651_d0_G16_mul1_G256_inv0 | ~t659_dec_1_inp;
  wire clk117;
  assign clk117 = dec_72[7] & clk;

  always @(posedge clk117) begin
    q0_0_G4_mul2_G16_mul1_G256_inv0_reg117 <= b0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk118;
  assign clk118 = dec_72[7] & clk;

  always @(posedge clk118) begin
    q0_0_G4_mul2_G16_mul1_G256_inv0_reg118 <= d0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk119;
  assign clk119 = ~dec_72[7] & clk;

  always @(posedge clk119) begin
    q0_0_G4_mul2_G16_mul1_G256_inv0_reg119 <= t639_b0_G4_mul2_G16_mul1_G256_inv0;
  end

  wire clk120;
  assign clk120 = ~dec_72[7] & clk;

  always @(posedge clk120) begin
    q0_0_G4_mul2_G16_mul1_G256_inv0_reg120 <= t650_d0_G4_mul2_G16_mul1_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg121 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg122 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg123 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg124 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg125 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg126 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg127 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg128 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg129 <= c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg130 <= dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg131 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg132 <= dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg133 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg134 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg135 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg136 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg137 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg138 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg139 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg140 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg141 <= c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg142 <= ~t226_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg143 <= t227_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg144 <= ~t228_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg145 <= t229_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg146 <= t234_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg147 <= t236_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg148 <= t237_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg149 <= t238_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg150 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg151 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg152 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg153 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg154 <= ~dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg155 <= t244_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg156 <= ~t245_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg157 <= t246_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg158 <= c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg159 <= t251_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg160 <= t252_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg161 <= ~t253_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg162 <= c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg163 <= ~t259_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg164 <= ~t260_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg165 <= t261_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg166 <= t265_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg167 <= t267_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg168 <= t268_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg169 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg170 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg171 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg172 <= y_reg171;
  end


  always @(posedge clk) begin
    y_reg173 <= t273_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg174 <= ~t275_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg175 <= t276_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg176 <= ~t277_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg177 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg178 <= t281_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg179 <= ~t287_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg180 <= t288_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg181 <= c0_G16_inv0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg182 <= ~dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg183 <= y_reg182;
  end


  always @(posedge clk) begin
    y_reg184 <= t294_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg185 <= y_reg184;
  end


  always @(posedge clk) begin
    y_reg186 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg187 <= y_reg186;
  end


  always @(posedge clk) begin
    y_reg188 <= t297_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg189 <= y_reg188;
  end


  always @(posedge clk) begin
    y_reg190 <= ~t298_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg191 <= y_reg190;
  end


  always @(posedge clk) begin
    y_reg192 <= t299_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg193 <= y_reg192;
  end


  always @(posedge clk) begin
    y_reg194 <= ~t304_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg195 <= t306_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg196 <= t307_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg197 <= t308_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg198 <= ~p0_0_G4_mul4_G16_inv0_G256_inv0_reg58;
  end


  always @(posedge clk) begin
    y_reg199 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg200 <= y_reg199;
  end


  always @(posedge clk) begin
    y_reg201 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg202 <= y_reg201;
  end


  always @(posedge clk) begin
    y_reg203 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg204 <= y_reg203;
  end


  always @(posedge clk) begin
    y_reg205 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg206 <= y_reg205;
  end


  always @(posedge clk) begin
    y_reg207 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg208 <= y_reg207;
  end


  always @(posedge clk) begin
    y_reg209 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg210 <= y_reg209;
  end


  always @(posedge clk) begin
    y_reg211 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg212 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg213 <= p0_0_G4_mul4_G16_inv0_G256_inv0_reg56;
  end


  always @(posedge clk) begin
    y_reg214 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg215 <= y_reg214;
  end


  always @(posedge clk) begin
    y_reg216 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg217 <= y_reg216;
  end


  always @(posedge clk) begin
    y_reg218 <= t315_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg219 <= y_reg218;
  end


  always @(posedge clk) begin
    y_reg220 <= t316_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg221 <= y_reg220;
  end


  always @(posedge clk) begin
    y_reg222 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg223 <= y_reg222;
  end


  always @(posedge clk) begin
    y_reg224 <= t321_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg225 <= y_reg224;
  end


  always @(posedge clk) begin
    y_reg226 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg227 <= y_reg226;
  end


  always @(posedge clk) begin
    y_reg228 <= t324_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg229 <= y_reg228;
  end


  always @(posedge clk) begin
    y_reg230 <= ~t325_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg231 <= y_reg230;
  end


  always @(posedge clk) begin
    y_reg232 <= ~c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg233 <= ~t331_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg234 <= ~t332_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg235 <= t333_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg236 <= ~t337_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg237 <= t339_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg238 <= t340_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg239 <= ~e0_G4_mul4_G16_inv0_G256_inv0_reg62;
  end


  always @(posedge clk) begin
    y_reg240 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg241 <= y_reg240;
  end


  always @(posedge clk) begin
    y_reg242 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg243 <= e0_G4_mul4_G16_inv0_G256_inv0_reg60;
  end


  always @(posedge clk) begin
    y_reg244 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg245 <= y_reg244;
  end


  always @(posedge clk) begin
    y_reg246 <= y_reg245;
  end


  always @(posedge clk) begin
    y_reg247 <= c0_G16_inv0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg248 <= ~t346_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg249 <= y_reg248;
  end


  always @(posedge clk) begin
    y_reg250 <= t347_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg251 <= y_reg250;
  end


  always @(posedge clk) begin
    y_reg252 <= c0_G16_inv0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg253 <= ~t351_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg254 <= y_reg253;
  end


  always @(posedge clk) begin
    y_reg255 <= t352_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg256 <= y_reg255;
  end


  always @(posedge clk) begin
    y_reg257 <= ~t353_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg258 <= y_reg257;
  end


  always @(posedge clk) begin
    y_reg259 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg260 <= t357_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg261 <= ~t363_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg262 <= ~t364_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg263 <= ~q0_0_G4_mul4_G16_inv0_G256_inv0_reg66;
  end


  always @(posedge clk) begin
    y_reg264 <= q0_0_G4_mul4_G16_inv0_G256_inv0_reg64;
  end


  always @(posedge clk) begin
    y_reg265 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg266 <= y_reg265;
  end


  always @(posedge clk) begin
    y_reg267 <= y_reg266;
  end


  always @(posedge clk) begin
    y_reg268 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg269 <= y_reg268;
  end


  always @(posedge clk) begin
    y_reg270 <= t370_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg271 <= y_reg270;
  end


  always @(posedge clk) begin
    y_reg272 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg273 <= y_reg272;
  end


  always @(posedge clk) begin
    y_reg274 <= t373_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg275 <= y_reg274;
  end


  always @(posedge clk) begin
    y_reg276 <= ~t374_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg277 <= y_reg276;
  end


  always @(posedge clk) begin
    y_reg278 <= t375_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg279 <= y_reg278;
  end


  always @(posedge clk) begin
    y_reg280 <= c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg281 <= t381_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg282 <= t382_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg283 <= ~t383_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg284 <= t384_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg285 <= ~p0_0_G4_mul5_G16_inv0_G256_inv0_reg70;
  end


  always @(posedge clk) begin
    y_reg286 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg287 <= y_reg286;
  end


  always @(posedge clk) begin
    y_reg288 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg289 <= y_reg288;
  end


  always @(posedge clk) begin
    y_reg290 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg291 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg292 <= p0_0_G4_mul5_G16_inv0_G256_inv0_reg68;
  end


  always @(posedge clk) begin
    y_reg293 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg294 <= y_reg293;
  end


  always @(posedge clk) begin
    y_reg295 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg296 <= y_reg295;
  end


  always @(posedge clk) begin
    y_reg297 <= t391_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg298 <= y_reg297;
  end


  always @(posedge clk) begin
    y_reg299 <= t392_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg300 <= y_reg299;
  end


  always @(posedge clk) begin
    y_reg301 <= ~dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg302 <= y_reg301;
  end


  always @(posedge clk) begin
    y_reg303 <= t397_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg304 <= y_reg303;
  end


  always @(posedge clk) begin
    y_reg305 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg306 <= y_reg305;
  end


  always @(posedge clk) begin
    y_reg307 <= t400_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg308 <= y_reg307;
  end


  always @(posedge clk) begin
    y_reg309 <= ~t401_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg310 <= y_reg309;
  end


  always @(posedge clk) begin
    y_reg311 <= dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg312 <= t407_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg313 <= t408_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg314 <= t409_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg315 <= ~c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg316 <= t414_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg317 <= t415_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg318 <= t416_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg319 <= ~e0_G4_mul5_G16_inv0_G256_inv0_reg76;
  end


  always @(posedge clk) begin
    y_reg320 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg321 <= y_reg320;
  end


  always @(posedge clk) begin
    y_reg322 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg323 <= cxord_0_G4_mul5_G16_inv0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg324 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg325 <= y_reg324;
  end


  always @(posedge clk) begin
    y_reg326 <= y_reg325;
  end


  always @(posedge clk) begin
    y_reg327 <= c0_G16_inv0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg328 <= ~t422_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg329 <= y_reg328;
  end


  always @(posedge clk) begin
    y_reg330 <= t423_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg331 <= y_reg330;
  end


  always @(posedge clk) begin
    y_reg332 <= c0_G16_inv0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg333 <= ~t427_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg334 <= y_reg333;
  end


  always @(posedge clk) begin
    y_reg335 <= t428_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg336 <= y_reg335;
  end


  always @(posedge clk) begin
    y_reg337 <= t429_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg338 <= y_reg337;
  end


  always @(posedge clk) begin
    y_reg339 <= t434_c0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg340 <= ~t436_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg341 <= t437_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg342 <= t438_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg343 <= ~q0_0_G4_mul5_G16_inv0_G256_inv0_reg80;
  end


  always @(posedge clk) begin
    y_reg344 <= q0_0_G4_mul5_G16_inv0_G256_inv0_reg78;
  end


  always @(posedge clk) begin
    y_reg345 <= t527_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg346 <= y_reg345;
  end


  always @(posedge clk) begin
    y_reg347 <= y_reg346;
  end


  always @(posedge clk) begin
    y_reg348 <= t528_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg349 <= y_reg348;
  end


  always @(posedge clk) begin
    y_reg350 <= y_reg349;
  end


  always @(posedge clk) begin
    y_reg351 <= t529_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg352 <= y_reg351;
  end


  always @(posedge clk) begin
    y_reg353 <= y_reg352;
  end


  always @(posedge clk) begin
    y_reg354 <= t530_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg355 <= y_reg354;
  end


  always @(posedge clk) begin
    y_reg356 <= y_reg355;
  end


  always @(posedge clk) begin
    y_reg357 <= ~p0_0_G4_mul1_G16_mul1_G256_inv0_reg98;
  end


  always @(posedge clk) begin
    y_reg358 <= y_reg357;
  end


  always @(posedge clk) begin
    y_reg359 <= y_reg358;
  end


  always @(posedge clk) begin
    y_reg360 <= dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg361 <= y_reg360;
  end


  always @(posedge clk) begin
    y_reg362 <= y_reg361;
  end


  always @(posedge clk) begin
    y_reg363 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg364 <= y_reg363;
  end


  always @(posedge clk) begin
    y_reg365 <= y_reg364;
  end


  always @(posedge clk) begin
    y_reg366 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg367 <= y_reg366;
  end


  always @(posedge clk) begin
    y_reg368 <= y_reg367;
  end


  always @(posedge clk) begin
    y_reg369 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg370 <= y_reg369;
  end


  always @(posedge clk) begin
    y_reg371 <= y_reg370;
  end


  always @(posedge clk) begin
    y_reg372 <= p0_0_G4_mul1_G16_mul1_G256_inv0_reg96;
  end


  always @(posedge clk) begin
    y_reg373 <= y_reg372;
  end


  always @(posedge clk) begin
    y_reg374 <= y_reg373;
  end


  always @(posedge clk) begin
    y_reg375 <= ~dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg376 <= y_reg375;
  end


  always @(posedge clk) begin
    y_reg377 <= y_reg376;
  end


  always @(posedge clk) begin
    y_reg378 <= t545_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg379 <= y_reg378;
  end


  always @(posedge clk) begin
    y_reg380 <= y_reg379;
  end


  always @(posedge clk) begin
    y_reg381 <= ~t546_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg382 <= y_reg381;
  end


  always @(posedge clk) begin
    y_reg383 <= y_reg382;
  end


  always @(posedge clk) begin
    y_reg384 <= t547_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg385 <= y_reg384;
  end


  always @(posedge clk) begin
    y_reg386 <= y_reg385;
  end


  always @(posedge clk) begin
    y_reg387 <= ~t552_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg388 <= y_reg387;
  end


  always @(posedge clk) begin
    y_reg389 <= y_reg388;
  end


  always @(posedge clk) begin
    y_reg390 <= t553_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg391 <= y_reg390;
  end


  always @(posedge clk) begin
    y_reg392 <= y_reg391;
  end


  always @(posedge clk) begin
    y_reg393 <= ~t554_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg394 <= y_reg393;
  end


  always @(posedge clk) begin
    y_reg395 <= y_reg394;
  end


  always @(posedge clk) begin
    y_reg396 <= ~e0_G4_mul1_G16_mul1_G256_inv0_reg104;
  end


  always @(posedge clk) begin
    y_reg397 <= y_reg396;
  end


  always @(posedge clk) begin
    y_reg398 <= y_reg397;
  end


  always @(posedge clk) begin
    y_reg399 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg400 <= y_reg399;
  end


  always @(posedge clk) begin
    y_reg401 <= y_reg400;
  end


  always @(posedge clk) begin
    y_reg402 <= cxord_0_G4_mul1_G16_mul1_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg403 <= y_reg402;
  end


  always @(posedge clk) begin
    y_reg404 <= y_reg403;
  end


  always @(posedge clk) begin
    y_reg405 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg406 <= y_reg405;
  end


  always @(posedge clk) begin
    y_reg407 <= y_reg406;
  end


  always @(posedge clk) begin
    y_reg408 <= y_reg407;
  end


  always @(posedge clk) begin
    y_reg409 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg410 <= y_reg409;
  end


  always @(posedge clk) begin
    y_reg411 <= y_reg410;
  end


  always @(posedge clk) begin
    y_reg412 <= ~t576_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg413 <= y_reg412;
  end


  always @(posedge clk) begin
    y_reg414 <= y_reg413;
  end


  always @(posedge clk) begin
    y_reg415 <= t577_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg416 <= y_reg415;
  end


  always @(posedge clk) begin
    y_reg417 <= y_reg416;
  end


  always @(posedge clk) begin
    y_reg418 <= ~t578_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg419 <= y_reg418;
  end


  always @(posedge clk) begin
    y_reg420 <= y_reg419;
  end


  always @(posedge clk) begin
    y_reg421 <= ~q0_0_G4_mul1_G16_mul1_G256_inv0_reg108;
  end


  always @(posedge clk) begin
    y_reg422 <= y_reg421;
  end


  always @(posedge clk) begin
    y_reg423 <= y_reg422;
  end


  always @(posedge clk) begin
    y_reg424 <= q0_0_G4_mul1_G16_mul1_G256_inv0_reg106;
  end


  always @(posedge clk) begin
    y_reg425 <= y_reg424;
  end


  always @(posedge clk) begin
    y_reg426 <= y_reg425;
  end


  always @(posedge clk) begin
    y_reg427 <= ~dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg428 <= y_reg427;
  end


  always @(posedge clk) begin
    y_reg429 <= y_reg428;
  end


  always @(posedge clk) begin
    y_reg430 <= t444_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg431 <= y_reg430;
  end


  always @(posedge clk) begin
    y_reg432 <= y_reg431;
  end


  always @(posedge clk) begin
    y_reg433 <= t447_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg434 <= y_reg433;
  end


  always @(posedge clk) begin
    y_reg435 <= y_reg434;
  end


  always @(posedge clk) begin
    y_reg436 <= ~t448_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg437 <= y_reg436;
  end


  always @(posedge clk) begin
    y_reg438 <= y_reg437;
  end


  always @(posedge clk) begin
    y_reg439 <= t449_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg440 <= y_reg439;
  end


  always @(posedge clk) begin
    y_reg441 <= y_reg440;
  end


  always @(posedge clk) begin
    y_reg442 <= ~p0_0_G4_mul0_G16_mul1_G256_inv0_reg84;
  end


  always @(posedge clk) begin
    y_reg443 <= y_reg442;
  end


  always @(posedge clk) begin
    y_reg444 <= y_reg443;
  end


  always @(posedge clk) begin
    y_reg445 <= dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg446 <= y_reg445;
  end


  always @(posedge clk) begin
    y_reg447 <= y_reg446;
  end


  always @(posedge clk) begin
    y_reg448 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg449 <= y_reg448;
  end


  always @(posedge clk) begin
    y_reg450 <= y_reg449;
  end


  always @(posedge clk) begin
    y_reg451 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg452 <= y_reg451;
  end


  always @(posedge clk) begin
    y_reg453 <= y_reg452;
  end


  always @(posedge clk) begin
    y_reg454 <= p0_0_G4_mul0_G16_mul1_G256_inv0_reg82;
  end


  always @(posedge clk) begin
    y_reg455 <= y_reg454;
  end


  always @(posedge clk) begin
    y_reg456 <= y_reg455;
  end


  always @(posedge clk) begin
    y_reg457 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg458 <= y_reg457;
  end


  always @(posedge clk) begin
    y_reg459 <= y_reg458;
  end


  always @(posedge clk) begin
    y_reg460 <= dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg461 <= y_reg460;
  end


  always @(posedge clk) begin
    y_reg462 <= y_reg461;
  end


  always @(posedge clk) begin
    y_reg463 <= t467_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg464 <= y_reg463;
  end


  always @(posedge clk) begin
    y_reg465 <= y_reg464;
  end


  always @(posedge clk) begin
    y_reg466 <= t468_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg467 <= y_reg466;
  end


  always @(posedge clk) begin
    y_reg468 <= y_reg467;
  end


  always @(posedge clk) begin
    y_reg469 <= ~dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg470 <= y_reg469;
  end


  always @(posedge clk) begin
    y_reg471 <= y_reg470;
  end


  always @(posedge clk) begin
    y_reg472 <= t473_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg473 <= y_reg472;
  end


  always @(posedge clk) begin
    y_reg474 <= y_reg473;
  end


  always @(posedge clk) begin
    y_reg475 <= t476_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg476 <= y_reg475;
  end


  always @(posedge clk) begin
    y_reg477 <= y_reg476;
  end


  always @(posedge clk) begin
    y_reg478 <= ~t477_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg479 <= y_reg478;
  end


  always @(posedge clk) begin
    y_reg480 <= y_reg479;
  end


  always @(posedge clk) begin
    y_reg481 <= ~e0_G4_mul0_G16_mul1_G256_inv0_reg90;
  end


  always @(posedge clk) begin
    y_reg482 <= y_reg481;
  end


  always @(posedge clk) begin
    y_reg483 <= y_reg482;
  end


  always @(posedge clk) begin
    y_reg484 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg485 <= y_reg484;
  end


  always @(posedge clk) begin
    y_reg486 <= y_reg485;
  end


  always @(posedge clk) begin
    y_reg487 <= cxord_0_G4_mul0_G16_mul1_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg488 <= y_reg487;
  end


  always @(posedge clk) begin
    y_reg489 <= y_reg488;
  end


  always @(posedge clk) begin
    y_reg490 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg491 <= y_reg490;
  end


  always @(posedge clk) begin
    y_reg492 <= y_reg491;
  end


  always @(posedge clk) begin
    y_reg493 <= y_reg492;
  end


  always @(posedge clk) begin
    y_reg494 <= t500_dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg495 <= y_reg494;
  end


  always @(posedge clk) begin
    y_reg496 <= y_reg495;
  end


  always @(posedge clk) begin
    y_reg497 <= t501_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg498 <= y_reg497;
  end


  always @(posedge clk) begin
    y_reg499 <= y_reg498;
  end


  always @(posedge clk) begin
    y_reg500 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg501 <= y_reg500;
  end


  always @(posedge clk) begin
    y_reg502 <= y_reg501;
  end


  always @(posedge clk) begin
    y_reg503 <= ~t506_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg504 <= y_reg503;
  end


  always @(posedge clk) begin
    y_reg505 <= y_reg504;
  end


  always @(posedge clk) begin
    y_reg506 <= t507_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg507 <= y_reg506;
  end


  always @(posedge clk) begin
    y_reg508 <= y_reg507;
  end


  always @(posedge clk) begin
    y_reg509 <= q0_0_G4_mul0_G16_mul1_G256_inv0_reg94;
  end


  always @(posedge clk) begin
    y_reg510 <= y_reg509;
  end


  always @(posedge clk) begin
    y_reg511 <= y_reg510;
  end


  always @(posedge clk) begin
    y_reg512 <= q0_0_G4_mul0_G16_mul1_G256_inv0_reg92;
  end


  always @(posedge clk) begin
    y_reg513 <= y_reg512;
  end


  always @(posedge clk) begin
    y_reg514 <= y_reg513;
  end


  always @(posedge clk) begin
    y_reg515 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg516 <= y_reg515;
  end


  always @(posedge clk) begin
    y_reg517 <= y_reg516;
  end


  always @(posedge clk) begin
    y_reg518 <= y_reg517;
  end


  always @(posedge clk) begin
    y_reg519 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg520 <= y_reg519;
  end


  always @(posedge clk) begin
    y_reg521 <= y_reg520;
  end


  always @(posedge clk) begin
    y_reg522 <= y_reg521;
  end


  always @(posedge clk) begin
    y_reg523 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg524 <= y_reg523;
  end


  always @(posedge clk) begin
    y_reg525 <= y_reg524;
  end


  always @(posedge clk) begin
    y_reg526 <= y_reg525;
  end


  always @(posedge clk) begin
    y_reg527 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg528 <= y_reg527;
  end


  always @(posedge clk) begin
    y_reg529 <= y_reg528;
  end


  always @(posedge clk) begin
    y_reg530 <= y_reg529;
  end


  always @(posedge clk) begin
    y_reg531 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg532 <= y_reg531;
  end


  always @(posedge clk) begin
    y_reg533 <= y_reg532;
  end


  always @(posedge clk) begin
    y_reg534 <= y_reg533;
  end


  always @(posedge clk) begin
    y_reg535 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg536 <= y_reg535;
  end


  always @(posedge clk) begin
    y_reg537 <= y_reg536;
  end


  always @(posedge clk) begin
    y_reg538 <= ~t595_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg539 <= y_reg538;
  end


  always @(posedge clk) begin
    y_reg540 <= y_reg539;
  end


  always @(posedge clk) begin
    y_reg541 <= ~t596_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg542 <= y_reg541;
  end


  always @(posedge clk) begin
    y_reg543 <= y_reg542;
  end


  always @(posedge clk) begin
    y_reg544 <= t597_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg545 <= y_reg544;
  end


  always @(posedge clk) begin
    y_reg546 <= y_reg545;
  end


  always @(posedge clk) begin
    y_reg547 <= ~p0_0_G4_mul2_G16_mul1_G256_inv0_reg112;
  end


  always @(posedge clk) begin
    y_reg548 <= y_reg547;
  end


  always @(posedge clk) begin
    y_reg549 <= y_reg548;
  end


  always @(posedge clk) begin
    y_reg550 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg551 <= y_reg550;
  end


  always @(posedge clk) begin
    y_reg552 <= y_reg551;
  end


  always @(posedge clk) begin
    y_reg553 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg554 <= y_reg553;
  end


  always @(posedge clk) begin
    y_reg555 <= y_reg554;
  end


  always @(posedge clk) begin
    y_reg556 <= p0_0_G4_mul2_G16_mul1_G256_inv0_reg110;
  end


  always @(posedge clk) begin
    y_reg557 <= y_reg556;
  end


  always @(posedge clk) begin
    y_reg558 <= y_reg557;
  end


  always @(posedge clk) begin
    y_reg559 <= t613_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg560 <= y_reg559;
  end


  always @(posedge clk) begin
    y_reg561 <= y_reg560;
  end


  always @(posedge clk) begin
    y_reg562 <= ~t614_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg563 <= y_reg562;
  end


  always @(posedge clk) begin
    y_reg564 <= y_reg563;
  end


  always @(posedge clk) begin
    y_reg565 <= t615_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg566 <= y_reg565;
  end


  always @(posedge clk) begin
    y_reg567 <= y_reg566;
  end


  always @(posedge clk) begin
    y_reg568 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg569 <= y_reg568;
  end


  always @(posedge clk) begin
    y_reg570 <= y_reg569;
  end


  always @(posedge clk) begin
    y_reg571 <= ~t621_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg572 <= y_reg571;
  end


  always @(posedge clk) begin
    y_reg573 <= y_reg572;
  end


  always @(posedge clk) begin
    y_reg574 <= ~t622_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg575 <= y_reg574;
  end


  always @(posedge clk) begin
    y_reg576 <= y_reg575;
  end


  always @(posedge clk) begin
    y_reg577 <= ~e0_G4_mul2_G16_mul1_G256_inv0_reg116;
  end


  always @(posedge clk) begin
    y_reg578 <= y_reg577;
  end


  always @(posedge clk) begin
    y_reg579 <= y_reg578;
  end


  always @(posedge clk) begin
    y_reg580 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg581 <= y_reg580;
  end


  always @(posedge clk) begin
    y_reg582 <= y_reg581;
  end


  always @(posedge clk) begin
    y_reg583 <= e0_G4_mul2_G16_mul1_G256_inv0_reg114;
  end


  always @(posedge clk) begin
    y_reg584 <= y_reg583;
  end


  always @(posedge clk) begin
    y_reg585 <= y_reg584;
  end


  always @(posedge clk) begin
    y_reg586 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg587 <= y_reg586;
  end


  always @(posedge clk) begin
    y_reg588 <= y_reg587;
  end


  always @(posedge clk) begin
    y_reg589 <= y_reg588;
  end


  always @(posedge clk) begin
    y_reg590 <= t644_dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg591 <= y_reg590;
  end


  always @(posedge clk) begin
    y_reg592 <= y_reg591;
  end


  always @(posedge clk) begin
    y_reg593 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg594 <= y_reg593;
  end


  always @(posedge clk) begin
    y_reg595 <= y_reg594;
  end


  always @(posedge clk) begin
    y_reg596 <= t648_dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg597 <= y_reg596;
  end


  always @(posedge clk) begin
    y_reg598 <= y_reg597;
  end


  always @(posedge clk) begin
    y_reg599 <= ~t649_dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg600 <= y_reg599;
  end


  always @(posedge clk) begin
    y_reg601 <= y_reg600;
  end


  always @(posedge clk) begin
    y_reg602 <= ~q0_0_G4_mul2_G16_mul1_G256_inv0_reg120;
  end


  always @(posedge clk) begin
    y_reg603 <= y_reg602;
  end


  always @(posedge clk) begin
    y_reg604 <= y_reg603;
  end


  always @(posedge clk) begin
    y_reg605 <= q0_0_G4_mul2_G16_mul1_G256_inv0_reg118;
  end


  always @(posedge clk) begin
    y_reg606 <= y_reg605;
  end


  always @(posedge clk) begin
    y_reg607 <= y_reg606;
  end


  always @(posedge clk) begin
    y_reg608 <= dec_4_inp;
  end


  always @(posedge clk) begin
    y_reg609 <= y_reg608;
  end


  always @(posedge clk) begin
    y_reg610 <= y_reg609;
  end


  always @(posedge clk) begin
    y_reg611 <= y_reg610;
  end


  always @(posedge clk) begin
    y_reg612 <= dec_12_inp;
  end


  always @(posedge clk) begin
    y_reg613 <= y_reg612;
  end


  always @(posedge clk) begin
    y_reg614 <= y_reg613;
  end


  always @(posedge clk) begin
    y_reg615 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg616 <= y_reg615;
  end


  always @(posedge clk) begin
    y_reg617 <= y_reg616;
  end


  always @(posedge clk) begin
    y_reg618 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg619 <= y_reg618;
  end


  always @(posedge clk) begin
    y_reg620 <= y_reg619;
  end


  always @(posedge clk) begin
    y_reg621 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg622 <= y_reg621;
  end


  always @(posedge clk) begin
    y_reg623 <= y_reg622;
  end


  always @(posedge clk) begin
    y_reg624 <= c0_G4_mul1_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg625 <= y_reg624;
  end


  always @(posedge clk) begin
    y_reg626 <= y_reg625;
  end


  always @(posedge clk) begin
    y_reg627 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg628 <= y_reg627;
  end


  always @(posedge clk) begin
    y_reg629 <= y_reg628;
  end


  always @(posedge clk) begin
    y_reg630 <= cxord_0_G4_mul1_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg631 <= y_reg630;
  end


  always @(posedge clk) begin
    y_reg632 <= y_reg631;
  end


  always @(posedge clk) begin
    y_reg633 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg634 <= y_reg633;
  end


  always @(posedge clk) begin
    y_reg635 <= y_reg634;
  end


  always @(posedge clk) begin
    y_reg636 <= d0_G4_mul1_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg637 <= y_reg636;
  end


  always @(posedge clk) begin
    y_reg638 <= y_reg637;
  end


  always @(posedge clk) begin
    y_reg639 <= dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg640 <= y_reg639;
  end


  always @(posedge clk) begin
    y_reg641 <= y_reg640;
  end


  always @(posedge clk) begin
    y_reg642 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg643 <= y_reg642;
  end


  always @(posedge clk) begin
    y_reg644 <= y_reg643;
  end


  always @(posedge clk) begin
    y_reg645 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg646 <= y_reg645;
  end


  always @(posedge clk) begin
    y_reg647 <= y_reg646;
  end


  always @(posedge clk) begin
    y_reg648 <= c0_G4_mul0_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg649 <= y_reg648;
  end


  always @(posedge clk) begin
    y_reg650 <= y_reg649;
  end


  always @(posedge clk) begin
    y_reg651 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg652 <= y_reg651;
  end


  always @(posedge clk) begin
    y_reg653 <= y_reg652;
  end


  always @(posedge clk) begin
    y_reg654 <= cxord_0_G4_mul0_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg655 <= y_reg654;
  end


  always @(posedge clk) begin
    y_reg656 <= y_reg655;
  end


  always @(posedge clk) begin
    y_reg657 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg658 <= y_reg657;
  end


  always @(posedge clk) begin
    y_reg659 <= y_reg658;
  end


  always @(posedge clk) begin
    y_reg660 <= d0_G4_mul0_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg661 <= y_reg660;
  end


  always @(posedge clk) begin
    y_reg662 <= y_reg661;
  end


  always @(posedge clk) begin
    y_reg663 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg664 <= y_reg663;
  end


  always @(posedge clk) begin
    y_reg665 <= y_reg664;
  end


  always @(posedge clk) begin
    y_reg666 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg667 <= y_reg666;
  end


  always @(posedge clk) begin
    y_reg668 <= y_reg667;
  end


  always @(posedge clk) begin
    y_reg669 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg670 <= y_reg669;
  end


  always @(posedge clk) begin
    y_reg671 <= y_reg670;
  end


  always @(posedge clk) begin
    y_reg672 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg673 <= y_reg672;
  end


  always @(posedge clk) begin
    y_reg674 <= y_reg673;
  end


  always @(posedge clk) begin
    y_reg675 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg676 <= y_reg675;
  end


  always @(posedge clk) begin
    y_reg677 <= y_reg676;
  end


  always @(posedge clk) begin
    y_reg678 <= dec_2_inp;
  end


  always @(posedge clk) begin
    y_reg679 <= y_reg678;
  end


  always @(posedge clk) begin
    y_reg680 <= y_reg679;
  end


  always @(posedge clk) begin
    y_reg681 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg682 <= y_reg681;
  end


  always @(posedge clk) begin
    y_reg683 <= y_reg682;
  end


  always @(posedge clk) begin
    y_reg684 <= c0_G4_mul2_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg685 <= y_reg684;
  end


  always @(posedge clk) begin
    y_reg686 <= y_reg685;
  end


  always @(posedge clk) begin
    y_reg687 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg688 <= y_reg687;
  end


  always @(posedge clk) begin
    y_reg689 <= y_reg688;
  end


  always @(posedge clk) begin
    y_reg690 <= cxord_0_G4_mul2_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg691 <= y_reg690;
  end


  always @(posedge clk) begin
    y_reg692 <= y_reg691;
  end


  always @(posedge clk) begin
    y_reg693 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg694 <= y_reg693;
  end


  always @(posedge clk) begin
    y_reg695 <= y_reg694;
  end


  always @(posedge clk) begin
    y_reg696 <= d0_G4_mul2_G16_mul2_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg697 <= y_reg696;
  end


  always @(posedge clk) begin
    y_reg698 <= y_reg697;
  end


  always @(posedge clk) begin
    y_reg699 <= q0_G256_inv0;
  end


  always @(posedge clk) begin
    y_reg700 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg701 <= y_reg700;
  end


  always @(posedge clk) begin
    y_reg702 <= y_reg701;
  end


  always @(posedge clk) begin
    y_reg703 <= y_reg702;
  end


  always @(posedge clk) begin
    y_reg704 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg705 <= y_reg704;
  end


  always @(posedge clk) begin
    y_reg706 <= y_reg705;
  end


  always @(posedge clk) begin
    y_reg707 <= y_reg706;
  end


  always @(posedge clk) begin
    y_reg708 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg709 <= y_reg708;
  end


  always @(posedge clk) begin
    y_reg710 <= y_reg709;
  end


  always @(posedge clk) begin
    y_reg711 <= y_reg710;
  end


  always @(posedge clk) begin
    y_reg712 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg713 <= y_reg712;
  end


  always @(posedge clk) begin
    y_reg714 <= y_reg713;
  end


  always @(posedge clk) begin
    y_reg715 <= y_reg714;
  end


  always @(posedge clk) begin
    y_reg716 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg717 <= y_reg716;
  end


  always @(posedge clk) begin
    y_reg718 <= y_reg717;
  end


  always @(posedge clk) begin
    y_reg719 <= y_reg718;
  end


  always @(posedge clk) begin
    y_reg720 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg721 <= y_reg720;
  end


  always @(posedge clk) begin
    y_reg722 <= y_reg721;
  end


  always @(posedge clk) begin
    y_reg723 <= y_reg722;
  end


  always @(posedge clk) begin
    y_reg724 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg725 <= y_reg724;
  end


  always @(posedge clk) begin
    y_reg726 <= y_reg725;
  end


  always @(posedge clk) begin
    y_reg727 <= y_reg726;
  end


  always @(posedge clk) begin
    y_reg728 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg729 <= y_reg728;
  end


  always @(posedge clk) begin
    y_reg730 <= y_reg729;
  end


  always @(posedge clk) begin
    y_reg731 <= y_reg730;
  end


  always @(posedge clk) begin
    y_reg732 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg733 <= y_reg732;
  end


  always @(posedge clk) begin
    y_reg734 <= y_reg733;
  end


  always @(posedge clk) begin
    y_reg735 <= y_reg734;
  end


  always @(posedge clk) begin
    y_reg736 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg737 <= y_reg736;
  end


  always @(posedge clk) begin
    y_reg738 <= y_reg737;
  end


  always @(posedge clk) begin
    y_reg739 <= y_reg738;
  end


  always @(posedge clk) begin
    y_reg740 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg741 <= y_reg740;
  end


  always @(posedge clk) begin
    y_reg742 <= y_reg741;
  end


  always @(posedge clk) begin
    y_reg743 <= y_reg742;
  end


  always @(posedge clk) begin
    y_reg744 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg745 <= y_reg744;
  end


  always @(posedge clk) begin
    y_reg746 <= y_reg745;
  end


  always @(posedge clk) begin
    y_reg747 <= y_reg746;
  end


  always @(posedge clk) begin
    y_reg748 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg749 <= y_reg748;
  end


  always @(posedge clk) begin
    y_reg750 <= y_reg749;
  end


  always @(posedge clk) begin
    y_reg751 <= y_reg750;
  end


  always @(posedge clk) begin
    y_reg752 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg753 <= y_reg752;
  end


  always @(posedge clk) begin
    y_reg754 <= y_reg753;
  end


  always @(posedge clk) begin
    y_reg755 <= y_reg754;
  end


  always @(posedge clk) begin
    y_reg756 <= dec_1_inp;
  end


  always @(posedge clk) begin
    y_reg757 <= y_reg756;
  end


  always @(posedge clk) begin
    y_reg758 <= y_reg757;
  end


  always @(posedge clk) begin
    y_reg759 <= y_reg758;
  end


  always @(posedge clk) begin
    y_reg760 <= yxorb1_G256_newbasis1;
  end


  always @(posedge clk) begin
    y_reg761 <= y_reg760;
  end


  always @(posedge clk) begin
    y_reg762 <= y_reg761;
  end


  always @(posedge clk) begin
    y_reg763 <= y_reg762;
  end


  always @(posedge clk) begin
    y_reg764 <= tempy1_G256_newbasis1;
  end


  always @(posedge clk) begin
    y_reg765 <= y_reg764;
  end


  always @(posedge clk) begin
    y_reg766 <= y_reg765;
  end


  always @(posedge clk) begin
    y_reg767 <= y_reg766;
  end


  always @(posedge clk) begin
    y_reg768 <= dec_3_inp;
  end


  always @(posedge clk) begin
    y_reg769 <= y_reg768;
  end


  always @(posedge clk) begin
    y_reg770 <= y_reg769;
  end


  always @(posedge clk) begin
    y_reg771 <= y_reg770;
  end


  always @(posedge clk) begin
    y_reg772 <= dec_4_inp;
  end


  always @(posedge clk) begin
    y_reg773 <= y_reg772;
  end


  always @(posedge clk) begin
    y_reg774 <= y_reg773;
  end


  always @(posedge clk) begin
    y_reg775 <= y_reg774;
  end


  always @(posedge clk) begin
    y_reg776 <= dec_220_inp;
  end


  always @(posedge clk) begin
    y_reg777 <= y_reg776;
  end


  always @(posedge clk) begin
    y_reg778 <= y_reg777;
  end


  always @(posedge clk) begin
    y_reg779 <= y_reg778;
  end


  always @(posedge clk) begin
    y_reg780 <= dec_11_inp;
  end


  always @(posedge clk) begin
    y_reg781 <= y_reg780;
  end


  always @(posedge clk) begin
    y_reg782 <= y_reg781;
  end


  always @(posedge clk) begin
    y_reg783 <= y_reg782;
  end


  always @(posedge clk) begin
    y_reg784 <= dec_158_inp;
  end


  always @(posedge clk) begin
    y_reg785 <= y_reg784;
  end


  always @(posedge clk) begin
    y_reg786 <= y_reg785;
  end


  always @(posedge clk) begin
    y_reg787 <= y_reg786;
  end


  always @(posedge clk) begin
    y_reg788 <= dec_45_inp;
  end


  always @(posedge clk) begin
    y_reg789 <= y_reg788;
  end


  always @(posedge clk) begin
    y_reg790 <= y_reg789;
  end


  always @(posedge clk) begin
    y_reg791 <= y_reg790;
  end


  always @(posedge clk) begin
    y_reg792 <= dec_88_inp;
  end


  always @(posedge clk) begin
    y_reg793 <= y_reg792;
  end


  always @(posedge clk) begin
    y_reg794 <= y_reg793;
  end


  always @(posedge clk) begin
    y_reg795 <= y_reg794;
  end


  always @(posedge clk) begin
    y_reg796 <= dec_99_inp;
  end


  always @(posedge clk) begin
    y_reg797 <= y_reg796;
  end


  always @(posedge clk) begin
    y_reg798 <= y_reg797;
  end


  always @(posedge clk) begin
    y_reg799 <= y_reg798;
  end


endmodule


